magic
tech sky130A
magscale 1 2
timestamp 1753620013
<< obsli1 >>
rect 1104 2159 9108 9809
<< obsm1 >>
rect 14 2128 9738 9840
<< metal2 >>
rect 1306 11618 1362 12418
rect 4526 11618 4582 12418
rect 7102 11618 7158 12418
rect 9678 11618 9734 12418
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 8390 0 8446 800
<< obsm2 >>
rect 20 11562 1250 11778
rect 1418 11562 4470 11778
rect 4638 11562 7046 11778
rect 7214 11562 9622 11778
rect 20 856 9732 11562
rect 130 711 2538 856
rect 2706 711 5114 856
rect 5282 711 8334 856
rect 8502 711 9732 856
<< metal3 >>
rect 0 11568 800 11688
rect 9474 9528 10274 9648
rect 0 8848 800 8968
rect 9474 6808 10274 6928
rect 0 5448 800 5568
rect 9474 3408 10274 3528
rect 0 2728 800 2848
rect 9474 688 10274 808
<< obsm3 >>
rect 880 11488 9474 11658
rect 800 9728 9474 11488
rect 800 9448 9394 9728
rect 800 9048 9474 9448
rect 880 8768 9474 9048
rect 800 7008 9474 8768
rect 800 6728 9394 7008
rect 800 5648 9474 6728
rect 880 5368 9474 5648
rect 800 3608 9474 5368
rect 800 3328 9394 3608
rect 800 2928 9474 3328
rect 880 2648 9474 2928
rect 800 888 9474 2648
rect 800 715 9394 888
<< metal4 >>
rect 1944 2128 2264 9840
rect 2604 2128 2924 9840
rect 3944 2128 4264 9840
rect 4604 2128 4924 9840
rect 5944 2128 6264 9840
rect 6604 2128 6924 9840
rect 7944 2128 8264 9840
rect 8604 2128 8924 9840
<< metal5 >>
rect 1056 9340 9156 9660
rect 1056 8680 9156 9000
rect 1056 7436 9156 7756
rect 1056 6776 9156 7096
rect 1056 5532 9156 5852
rect 1056 4872 9156 5192
rect 1056 3628 9156 3948
rect 1056 2968 9156 3288
<< labels >>
rlabel metal4 s 2604 2128 2924 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4604 2128 4924 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 6604 2128 6924 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8604 2128 8924 9840 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3628 9156 3948 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5532 9156 5852 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 7436 9156 7756 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9340 9156 9660 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1944 2128 2264 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 3944 2128 4264 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 5944 2128 6264 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7944 2128 8264 9840 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2968 9156 3288 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4872 9156 5192 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 6776 9156 7096 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8680 9156 9000 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 9474 6808 10274 6928 6 a[0]
port 3 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 a[1]
port 4 nsew signal input
rlabel metal3 s 9474 9528 10274 9648 6 a[2]
port 5 nsew signal input
rlabel metal3 s 9474 688 10274 808 6 a[3]
port 6 nsew signal input
rlabel metal2 s 4526 11618 4582 12418 6 b[0]
port 7 nsew signal input
rlabel metal2 s 18 0 74 800 6 b[1]
port 8 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 b[2]
port 9 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 b[3]
port 10 nsew signal input
rlabel metal2 s 7102 11618 7158 12418 6 carry
port 11 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 out[0]
port 12 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 out[1]
port 13 nsew signal output
rlabel metal2 s 9678 11618 9734 12418 6 out[2]
port 14 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 out[3]
port 15 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 sel[0]
port 16 nsew signal input
rlabel metal2 s 1306 11618 1362 12418 6 sel[1]
port 17 nsew signal input
rlabel metal3 s 9474 3408 10274 3528 6 sel[2]
port 18 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 10274 12418
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 420438
string GDS_FILE /openlane/designs/alu/runs/RUN_2025.07.27_12.38.31/results/signoff/alu.magic.gds
string GDS_START 200546
<< end >>

