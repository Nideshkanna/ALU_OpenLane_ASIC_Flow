VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alu
  CLASS BLOCK ;
  FOREIGN alu ;
  ORIGIN 0.000 0.000 ;
  SIZE 51.370 BY 62.090 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.020 10.640 14.620 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.020 10.640 24.620 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.020 10.640 34.620 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.020 10.640 44.620 49.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 18.140 45.780 19.740 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 27.660 45.780 29.260 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 37.180 45.780 38.780 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 46.700 45.780 48.300 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.720 10.640 11.320 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.720 10.640 21.320 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.720 10.640 31.320 49.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.720 10.640 41.320 49.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 14.840 45.780 16.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 24.360 45.780 25.960 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 33.880 45.780 35.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 43.400 45.780 45.000 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.370 34.040 51.370 34.640 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.370 47.640 51.370 48.240 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.370 3.440 51.370 4.040 ;
    END
  END a[3]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 58.090 22.910 62.090 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END b[3]
  PIN carry
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 35.510 58.090 35.790 62.090 ;
    END
  END carry
  PIN out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END out[0]
  PIN out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 58.090 48.670 62.090 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END out[3]
  PIN sel[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END sel[0]
  PIN sel[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 6.530 58.090 6.810 62.090 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 47.370 17.040 51.370 17.640 ;
    END
  END sel[2]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 45.540 49.045 ;
      LAYER met1 ;
        RECT 0.070 10.640 48.690 49.200 ;
      LAYER met2 ;
        RECT 0.100 57.810 6.250 58.890 ;
        RECT 7.090 57.810 22.350 58.890 ;
        RECT 23.190 57.810 35.230 58.890 ;
        RECT 36.070 57.810 48.110 58.890 ;
        RECT 0.100 4.280 48.660 57.810 ;
        RECT 0.650 3.555 12.690 4.280 ;
        RECT 13.530 3.555 25.570 4.280 ;
        RECT 26.410 3.555 41.670 4.280 ;
        RECT 42.510 3.555 48.660 4.280 ;
      LAYER met3 ;
        RECT 4.400 57.440 47.370 58.290 ;
        RECT 4.000 48.640 47.370 57.440 ;
        RECT 4.000 47.240 46.970 48.640 ;
        RECT 4.000 45.240 47.370 47.240 ;
        RECT 4.400 43.840 47.370 45.240 ;
        RECT 4.000 35.040 47.370 43.840 ;
        RECT 4.000 33.640 46.970 35.040 ;
        RECT 4.000 28.240 47.370 33.640 ;
        RECT 4.400 26.840 47.370 28.240 ;
        RECT 4.000 18.040 47.370 26.840 ;
        RECT 4.000 16.640 46.970 18.040 ;
        RECT 4.000 14.640 47.370 16.640 ;
        RECT 4.400 13.240 47.370 14.640 ;
        RECT 4.000 4.440 47.370 13.240 ;
        RECT 4.000 3.575 46.970 4.440 ;
  END
END alu
END LIBRARY

