* NGSPICE file created from alu.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxtn_1 abstract view
.subckt sky130_fd_sc_hd__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt alu VGND VPWR a[0] a[1] a[2] a[3] b[0] b[1] b[2] b[3] carry out[0] out[1]
+ out[2] out[3] sel[0] sel[1] sel[2]
XFILLER_0_3_28 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_062_ _006_ _010_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_061_ _007_ _008_ _009_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_060_ net6 net2 VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput12 net12 VGND VGND VPWR VPWR carry sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_11 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_110_ _000_ _001_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dlxtn_1
XFILLER_0_1_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput13 net13 VGND VGND VPWR VPWR out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 net14 VGND VGND VPWR VPWR out[1] sky130_fd_sc_hd__clkbuf_4
X_099_ _037_ _038_ _044_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__a21o_1
Xoutput15 net15 VGND VGND VPWR VPWR out[2] sky130_fd_sc_hd__clkbuf_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_098_ _039_ _026_ _041_ _006_ _043_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput16 net16 VGND VGND VPWR VPWR out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_097_ _039_ _011_ _030_ _042_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_096_ _010_ _015_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__or2b_1
X_079_ _026_ _024_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__nor2_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_095_ _039_ _028_ _040_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__o21bai_1
X_078_ _023_ net10 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_094_ _023_ net10 net9 VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_077_ _023_ net10 _024_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__and3_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_093_ net7 net3 VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_076_ net5 net1 net10 net9 VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 a[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_059_ net5 net1 VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__nand2_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput2 a[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ _015_ _018_ _002_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__a21oi_1
X_058_ net6 net2 VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__xnor2_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_075_ net11 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__inv_2
Xinput3 a[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_1
X_091_ _015_ _018_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__or2_1
X_074_ _002_ _003_ _013_ _021_ _022_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__a32o_1
X_057_ net7 net3 VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_109_ _052_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_090_ _030_ _031_ _033_ _036_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__a211o_1
Xinput4 a[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_056_ net7 net3 VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__nand2_1
X_073_ net8 net4 VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__or2b_1
X_108_ net11 net10 VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 b[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_1
XFILLER_0_11_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_072_ _014_ _020_ _002_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a21oi_1
X_055_ net8 net4 VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_107_ _045_ _046_ _051_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__a21o_1
XFILLER_0_11_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_071_ _015_ _018_ _019_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__a21o_1
Xinput6 b[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_054_ net8 net4 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__or2_1
X_106_ _021_ _047_ _049_ _003_ _050_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__a221o_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_070_ net7 net3 VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__and2b_1
XTAP_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 b[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_1
Xinput10 sel[1] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_053_ net11 net10 net9 VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__or3b_2
X_105_ net8 net4 _026_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__and3_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 b[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XTAP_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput11 sel[2] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
X_104_ _040_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__or2_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 sel[0] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_11_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_103_ _028_ _004_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_102_ _014_ _020_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_101_ _014_ _012_ _030_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_100_ _014_ _012_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_089_ net6 net2 _026_ _034_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__o221a_1
XTAP_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ _023_ net10 _034_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_087_ net6 net2 net9 VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_086_ _007_ _016_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__o21ba_1
X_069_ _007_ _016_ _017_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_085_ _007_ _016_ _002_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__a21o_1
XFILLER_0_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_068_ net6 net2 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__and2b_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_067_ net1 net5 VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__or2b_1
XFILLER_0_9_22 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_084_ _007_ _008_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__xor2_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_083_ _002_ _028_ _029_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_066_ _005_ _006_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_065_ _004_ _003_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nand2_1
X_082_ _023_ net9 net10 VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_081_ _023_ net10 net9 VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__or3_1
XFILLER_0_10_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_064_ _004_ _012_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__nand2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_080_ net5 net1 _025_ _027_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__o22a_1
X_063_ _005_ _011_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
.ends

