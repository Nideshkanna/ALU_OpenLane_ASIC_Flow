magic
tech sky130A
magscale 1 2
timestamp 1753620023
<< checkpaint >>
rect -3932 -3932 14206 16350
<< viali >>
rect 1501 9605 1535 9639
rect 1869 9605 1903 9639
rect 7665 9605 7699 9639
rect 8401 9605 8435 9639
rect 8769 9605 8803 9639
rect 4629 9537 4663 9571
rect 7297 9537 7331 9571
rect 8217 9537 8251 9571
rect 1593 9333 1627 9367
rect 1961 9333 1995 9367
rect 4813 9333 4847 9367
rect 8033 9333 8067 9367
rect 6285 9129 6319 9163
rect 4997 9061 5031 9095
rect 5273 8993 5307 9027
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 3065 8925 3099 8959
rect 3341 8925 3375 8959
rect 3433 8925 3467 8959
rect 4077 8925 4111 8959
rect 4445 8925 4479 8959
rect 4813 8925 4847 8959
rect 5549 8925 5583 8959
rect 3249 8857 3283 8891
rect 4261 8857 4295 8891
rect 3617 8789 3651 8823
rect 3601 8585 3635 8619
rect 3801 8517 3835 8551
rect 2513 8449 2547 8483
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3065 8449 3099 8483
rect 3341 8449 3375 8483
rect 3985 8449 4019 8483
rect 4169 8449 4203 8483
rect 4721 8449 4755 8483
rect 2605 8381 2639 8415
rect 2789 8313 2823 8347
rect 3249 8313 3283 8347
rect 4077 8313 4111 8347
rect 3433 8245 3467 8279
rect 3617 8245 3651 8279
rect 4997 8245 5031 8279
rect 5181 8245 5215 8279
rect 7205 8041 7239 8075
rect 6377 7973 6411 8007
rect 1685 7905 1719 7939
rect 7665 7905 7699 7939
rect 1869 7837 1903 7871
rect 4813 7837 4847 7871
rect 5089 7837 5123 7871
rect 5365 7837 5399 7871
rect 5641 7837 5675 7871
rect 6653 7837 6687 7871
rect 6745 7837 6779 7871
rect 6837 7837 6871 7871
rect 7021 7837 7055 7871
rect 5273 7769 5307 7803
rect 6377 7769 6411 7803
rect 7297 7769 7331 7803
rect 7481 7769 7515 7803
rect 2513 7701 2547 7735
rect 4905 7701 4939 7735
rect 5457 7701 5491 7735
rect 5825 7701 5859 7735
rect 6561 7701 6595 7735
rect 3065 7497 3099 7531
rect 2605 7429 2639 7463
rect 6745 7429 6779 7463
rect 4813 7361 4847 7395
rect 5089 7361 5123 7395
rect 5273 7361 5307 7395
rect 6561 7361 6595 7395
rect 6837 7361 6871 7395
rect 8769 7361 8803 7395
rect 2881 7225 2915 7259
rect 8585 7225 8619 7259
rect 4629 7157 4663 7191
rect 6377 7157 6411 7191
rect 7941 6953 7975 6987
rect 8033 6885 8067 6919
rect 8401 6681 8435 6715
rect 1777 6409 1811 6443
rect 2789 6409 2823 6443
rect 7389 6409 7423 6443
rect 8309 6341 8343 6375
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 2053 6273 2087 6307
rect 2241 6273 2275 6307
rect 2605 6273 2639 6307
rect 2881 6273 2915 6307
rect 3065 6273 3099 6307
rect 3617 6273 3651 6307
rect 4261 6273 4295 6307
rect 4353 6273 4387 6307
rect 4537 6273 4571 6307
rect 4629 6273 4663 6307
rect 4997 6273 5031 6307
rect 6101 6273 6135 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 7389 6273 7423 6307
rect 7573 6273 7607 6307
rect 8125 6273 8159 6307
rect 2329 6205 2363 6239
rect 2421 6205 2455 6239
rect 3709 6205 3743 6239
rect 3985 6205 4019 6239
rect 4721 6205 4755 6239
rect 7941 6205 7975 6239
rect 1961 6137 1995 6171
rect 2973 6137 3007 6171
rect 4813 6137 4847 6171
rect 4077 6069 4111 6103
rect 4905 6069 4939 6103
rect 5641 6069 5675 6103
rect 5825 6069 5859 6103
rect 6469 6069 6503 6103
rect 1777 5865 1811 5899
rect 6745 5865 6779 5899
rect 7941 5865 7975 5899
rect 8493 5797 8527 5831
rect 1961 5729 1995 5763
rect 7757 5729 7791 5763
rect 1685 5661 1719 5695
rect 5365 5661 5399 5695
rect 5549 5661 5583 5695
rect 5641 5661 5675 5695
rect 5733 5661 5767 5695
rect 6101 5661 6135 5695
rect 6249 5661 6283 5695
rect 6469 5661 6503 5695
rect 6566 5661 6600 5695
rect 7573 5661 7607 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 8401 5661 8435 5695
rect 8585 5661 8619 5695
rect 6009 5593 6043 5627
rect 6377 5593 6411 5627
rect 1961 5525 1995 5559
rect 7389 5525 7423 5559
rect 3157 5321 3191 5355
rect 4997 5321 5031 5355
rect 1409 5253 1443 5287
rect 1777 5253 1811 5287
rect 3249 5185 3283 5219
rect 5089 5185 5123 5219
rect 5273 5185 5307 5219
rect 4813 4981 4847 5015
rect 2329 4777 2363 4811
rect 2973 4777 3007 4811
rect 3433 4777 3467 4811
rect 3617 4777 3651 4811
rect 3985 4777 4019 4811
rect 3157 4709 3191 4743
rect 4629 4709 4663 4743
rect 4813 4709 4847 4743
rect 2513 4641 2547 4675
rect 4353 4641 4387 4675
rect 1869 4573 1903 4607
rect 1961 4573 1995 4607
rect 2237 4573 2271 4607
rect 3249 4573 3283 4607
rect 3341 4573 3375 4607
rect 5089 4573 5123 4607
rect 3019 4539 3053 4573
rect 2789 4505 2823 4539
rect 3801 4505 3835 4539
rect 4905 4505 4939 4539
rect 2145 4437 2179 4471
rect 2513 4437 2547 4471
rect 4001 4437 4035 4471
rect 4169 4437 4203 4471
rect 5273 4437 5307 4471
rect 3249 4233 3283 4267
rect 5917 4165 5951 4199
rect 6377 4165 6411 4199
rect 3065 4097 3099 4131
rect 5339 4097 5373 4131
rect 5457 4097 5491 4131
rect 5549 4097 5583 4131
rect 5641 4097 5675 4131
rect 6101 4097 6135 4131
rect 6193 4097 6227 4131
rect 6561 4097 6595 4131
rect 7205 4097 7239 4131
rect 7389 4097 7423 4131
rect 7573 4097 7607 4131
rect 7757 4097 7791 4131
rect 3433 4029 3467 4063
rect 5181 4029 5215 4063
rect 7481 4029 7515 4063
rect 5917 3961 5951 3995
rect 7665 3961 7699 3995
rect 3433 3893 3467 3927
rect 5825 3893 5859 3927
rect 6745 3893 6779 3927
rect 7021 3893 7055 3927
rect 8585 3621 8619 3655
rect 5641 3485 5675 3519
rect 5734 3485 5768 3519
rect 6147 3485 6181 3519
rect 8769 3485 8803 3519
rect 5917 3417 5951 3451
rect 6009 3417 6043 3451
rect 6285 3349 6319 3383
rect 4169 3145 4203 3179
rect 4905 3145 4939 3179
rect 5197 3145 5231 3179
rect 5365 3145 5399 3179
rect 5825 3145 5859 3179
rect 6193 3145 6227 3179
rect 1777 3077 1811 3111
rect 4997 3077 5031 3111
rect 4169 3009 4203 3043
rect 4353 3009 4387 3043
rect 4445 3009 4479 3043
rect 5457 3009 5491 3043
rect 5641 3009 5675 3043
rect 6009 3009 6043 3043
rect 6193 3009 6227 3043
rect 6653 3009 6687 3043
rect 6837 3009 6871 3043
rect 6929 3009 6963 3043
rect 7205 3009 7239 3043
rect 7389 3009 7423 3043
rect 7297 2941 7331 2975
rect 1501 2805 1535 2839
rect 4537 2805 4571 2839
rect 5181 2805 5215 2839
rect 6469 2805 6503 2839
rect 1593 2601 1627 2635
rect 2881 2601 2915 2635
rect 8217 2601 8251 2635
rect 8677 2601 8711 2635
rect 2697 2397 2731 2431
rect 5457 2397 5491 2431
rect 8401 2397 8435 2431
rect 8493 2397 8527 2431
rect 1501 2329 1535 2363
rect 5181 2261 5215 2295
<< metal1 >>
rect 1104 9818 9108 9840
rect 1104 9766 2610 9818
rect 2662 9766 2674 9818
rect 2726 9766 2738 9818
rect 2790 9766 2802 9818
rect 2854 9766 2866 9818
rect 2918 9766 4610 9818
rect 4662 9766 4674 9818
rect 4726 9766 4738 9818
rect 4790 9766 4802 9818
rect 4854 9766 4866 9818
rect 4918 9766 6610 9818
rect 6662 9766 6674 9818
rect 6726 9766 6738 9818
rect 6790 9766 6802 9818
rect 6854 9766 6866 9818
rect 6918 9766 8610 9818
rect 8662 9766 8674 9818
rect 8726 9766 8738 9818
rect 8790 9766 8802 9818
rect 8854 9766 8866 9818
rect 8918 9766 9108 9818
rect 1104 9744 9108 9766
rect 1302 9596 1308 9648
rect 1360 9636 1366 9648
rect 1489 9639 1547 9645
rect 1489 9636 1501 9639
rect 1360 9608 1501 9636
rect 1360 9596 1366 9608
rect 1489 9605 1501 9608
rect 1535 9605 1547 9639
rect 1489 9599 1547 9605
rect 1854 9596 1860 9648
rect 1912 9596 1918 9648
rect 4522 9596 4528 9648
rect 4580 9596 4586 9648
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 7653 9639 7711 9645
rect 7653 9636 7665 9639
rect 7432 9608 7665 9636
rect 7432 9596 7438 9608
rect 7653 9605 7665 9608
rect 7699 9605 7711 9639
rect 7653 9599 7711 9605
rect 7742 9596 7748 9648
rect 7800 9636 7806 9648
rect 8389 9639 8447 9645
rect 8389 9636 8401 9639
rect 7800 9608 8401 9636
rect 7800 9596 7806 9608
rect 8389 9605 8401 9608
rect 8435 9605 8447 9639
rect 8389 9599 8447 9605
rect 8757 9639 8815 9645
rect 8757 9605 8769 9639
rect 8803 9636 8815 9639
rect 9674 9636 9680 9648
rect 8803 9608 9680 9636
rect 8803 9605 8815 9608
rect 8757 9599 8815 9605
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 4540 9568 4568 9596
rect 4617 9571 4675 9577
rect 4617 9568 4629 9571
rect 4540 9540 4629 9568
rect 4617 9537 4629 9540
rect 4663 9537 4675 9571
rect 4617 9531 4675 9537
rect 7282 9528 7288 9580
rect 7340 9528 7346 9580
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9537 8263 9571
rect 8205 9531 8263 9537
rect 8220 9500 8248 9531
rect 8938 9528 8944 9580
rect 8996 9528 9002 9580
rect 8956 9500 8984 9528
rect 8220 9472 8984 9500
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1544 9336 1593 9364
rect 1544 9324 1550 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 1949 9367 2007 9373
rect 1949 9364 1961 9367
rect 1728 9336 1961 9364
rect 1728 9324 1734 9336
rect 1949 9333 1961 9336
rect 1995 9333 2007 9367
rect 1949 9327 2007 9333
rect 4801 9367 4859 9373
rect 4801 9333 4813 9367
rect 4847 9364 4859 9367
rect 4982 9364 4988 9376
rect 4847 9336 4988 9364
rect 4847 9333 4859 9336
rect 4801 9327 4859 9333
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 8021 9367 8079 9373
rect 8021 9364 8033 9367
rect 7892 9336 8033 9364
rect 7892 9324 7898 9336
rect 8021 9333 8033 9336
rect 8067 9333 8079 9367
rect 8021 9327 8079 9333
rect 1104 9274 9108 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 3950 9274
rect 4002 9222 4014 9274
rect 4066 9222 4078 9274
rect 4130 9222 4142 9274
rect 4194 9222 4206 9274
rect 4258 9222 5950 9274
rect 6002 9222 6014 9274
rect 6066 9222 6078 9274
rect 6130 9222 6142 9274
rect 6194 9222 6206 9274
rect 6258 9222 7950 9274
rect 8002 9222 8014 9274
rect 8066 9222 8078 9274
rect 8130 9222 8142 9274
rect 8194 9222 8206 9274
rect 8258 9222 9108 9274
rect 1104 9200 9108 9222
rect 6273 9163 6331 9169
rect 6273 9129 6285 9163
rect 6319 9160 6331 9163
rect 7282 9160 7288 9172
rect 6319 9132 7288 9160
rect 6319 9129 6331 9132
rect 6273 9123 6331 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 4985 9095 5043 9101
rect 4985 9061 4997 9095
rect 5031 9061 5043 9095
rect 4985 9055 5043 9061
rect 3510 9024 3516 9036
rect 3252 8996 3516 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 1762 8956 1768 8968
rect 1719 8928 1768 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 1762 8916 1768 8928
rect 1820 8956 1826 8968
rect 3053 8959 3111 8965
rect 3053 8956 3065 8959
rect 1820 8928 3065 8956
rect 1820 8916 1826 8928
rect 3053 8925 3065 8928
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 1486 8848 1492 8900
rect 1544 8888 1550 8900
rect 3252 8897 3280 8996
rect 3510 8984 3516 8996
rect 3568 9024 3574 9036
rect 5000 9024 5028 9055
rect 5261 9027 5319 9033
rect 5261 9024 5273 9027
rect 3568 8996 4108 9024
rect 5000 8996 5273 9024
rect 3568 8984 3574 8996
rect 4080 8965 4108 8996
rect 5261 8993 5273 8996
rect 5307 8993 5319 9027
rect 5261 8987 5319 8993
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3421 8959 3479 8965
rect 3421 8925 3433 8959
rect 3467 8925 3479 8959
rect 3421 8919 3479 8925
rect 4065 8959 4123 8965
rect 4065 8925 4077 8959
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 3237 8891 3295 8897
rect 3237 8888 3249 8891
rect 1544 8860 3249 8888
rect 1544 8848 1550 8860
rect 3237 8857 3249 8860
rect 3283 8857 3295 8891
rect 3237 8851 3295 8857
rect 3344 8832 3372 8919
rect 3436 8888 3464 8919
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8956 4491 8959
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 4479 8928 4813 8956
rect 4479 8925 4491 8928
rect 4433 8919 4491 8925
rect 4801 8925 4813 8928
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8956 5595 8959
rect 5718 8956 5724 8968
rect 5583 8928 5724 8956
rect 5583 8925 5595 8928
rect 5537 8919 5595 8925
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 4172 8888 4200 8916
rect 3436 8860 4200 8888
rect 4249 8891 4307 8897
rect 4249 8857 4261 8891
rect 4295 8857 4307 8891
rect 4249 8851 4307 8857
rect 3326 8780 3332 8832
rect 3384 8780 3390 8832
rect 3418 8780 3424 8832
rect 3476 8820 3482 8832
rect 3602 8820 3608 8832
rect 3476 8792 3608 8820
rect 3476 8780 3482 8792
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 3694 8780 3700 8832
rect 3752 8820 3758 8832
rect 4264 8820 4292 8851
rect 3752 8792 4292 8820
rect 3752 8780 3758 8792
rect 1104 8730 9108 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 4610 8730
rect 4662 8678 4674 8730
rect 4726 8678 4738 8730
rect 4790 8678 4802 8730
rect 4854 8678 4866 8730
rect 4918 8678 6610 8730
rect 6662 8678 6674 8730
rect 6726 8678 6738 8730
rect 6790 8678 6802 8730
rect 6854 8678 6866 8730
rect 6918 8678 8610 8730
rect 8662 8678 8674 8730
rect 8726 8678 8738 8730
rect 8790 8678 8802 8730
rect 8854 8678 8866 8730
rect 8918 8678 9108 8730
rect 1104 8656 9108 8678
rect 3234 8616 3240 8628
rect 2700 8588 3240 8616
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 2700 8489 2728 8588
rect 3234 8576 3240 8588
rect 3292 8576 3298 8628
rect 3602 8625 3608 8628
rect 3589 8619 3608 8625
rect 3589 8585 3601 8619
rect 3589 8579 3608 8585
rect 3602 8576 3608 8579
rect 3660 8576 3666 8628
rect 4982 8576 4988 8628
rect 5040 8576 5046 8628
rect 3786 8508 3792 8560
rect 3844 8508 3850 8560
rect 3988 8520 4752 8548
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 2958 8440 2964 8492
rect 3016 8440 3022 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 2593 8415 2651 8421
rect 2593 8381 2605 8415
rect 2639 8412 2651 8415
rect 3068 8412 3096 8443
rect 3326 8440 3332 8492
rect 3384 8480 3390 8492
rect 3988 8489 4016 8520
rect 3973 8483 4031 8489
rect 3973 8480 3985 8483
rect 3384 8452 3985 8480
rect 3384 8440 3390 8452
rect 3973 8449 3985 8452
rect 4019 8449 4031 8483
rect 4154 8480 4160 8492
rect 3973 8443 4031 8449
rect 4080 8452 4160 8480
rect 4080 8412 4108 8452
rect 4154 8440 4160 8452
rect 4212 8480 4218 8492
rect 4724 8489 4752 8520
rect 4709 8483 4767 8489
rect 4212 8452 4660 8480
rect 4212 8440 4218 8452
rect 2639 8384 3096 8412
rect 3528 8384 4108 8412
rect 4632 8412 4660 8452
rect 4709 8449 4721 8483
rect 4755 8480 4767 8483
rect 5000 8480 5028 8576
rect 4755 8452 5028 8480
rect 4755 8449 4767 8452
rect 4709 8443 4767 8449
rect 4632 8384 5028 8412
rect 2639 8381 2651 8384
rect 2593 8375 2651 8381
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 3142 8344 3148 8356
rect 2823 8316 3148 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 3237 8347 3295 8353
rect 3237 8313 3249 8347
rect 3283 8344 3295 8347
rect 3528 8344 3556 8384
rect 3283 8316 3556 8344
rect 3283 8313 3295 8316
rect 3237 8307 3295 8313
rect 3694 8304 3700 8356
rect 3752 8344 3758 8356
rect 4065 8347 4123 8353
rect 4065 8344 4077 8347
rect 3752 8316 4077 8344
rect 3752 8304 3758 8316
rect 4065 8313 4077 8316
rect 4111 8313 4123 8347
rect 4065 8307 4123 8313
rect 5000 8288 5028 8384
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3421 8279 3479 8285
rect 3421 8276 3433 8279
rect 3016 8248 3433 8276
rect 3016 8236 3022 8248
rect 3421 8245 3433 8248
rect 3467 8245 3479 8279
rect 3421 8239 3479 8245
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 3605 8279 3663 8285
rect 3605 8276 3617 8279
rect 3568 8248 3617 8276
rect 3568 8236 3574 8248
rect 3605 8245 3617 8248
rect 3651 8245 3663 8279
rect 3605 8239 3663 8245
rect 4982 8236 4988 8288
rect 5040 8236 5046 8288
rect 5166 8236 5172 8288
rect 5224 8236 5230 8288
rect 1104 8186 9108 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 3950 8186
rect 4002 8134 4014 8186
rect 4066 8134 4078 8186
rect 4130 8134 4142 8186
rect 4194 8134 4206 8186
rect 4258 8134 5950 8186
rect 6002 8134 6014 8186
rect 6066 8134 6078 8186
rect 6130 8134 6142 8186
rect 6194 8134 6206 8186
rect 6258 8134 7950 8186
rect 8002 8134 8014 8186
rect 8066 8134 8078 8186
rect 8130 8134 8142 8186
rect 8194 8134 8206 8186
rect 8258 8134 9108 8186
rect 1104 8112 9108 8134
rect 7193 8075 7251 8081
rect 7193 8041 7205 8075
rect 7239 8072 7251 8075
rect 7742 8072 7748 8084
rect 7239 8044 7748 8072
rect 7239 8041 7251 8044
rect 7193 8035 7251 8041
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 6365 8007 6423 8013
rect 6365 7973 6377 8007
rect 6411 7973 6423 8007
rect 6365 7967 6423 7973
rect 1670 7896 1676 7948
rect 1728 7896 1734 7948
rect 5166 7936 5172 7948
rect 4816 7908 5172 7936
rect 1854 7828 1860 7880
rect 1912 7828 1918 7880
rect 4816 7877 4844 7908
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 6380 7936 6408 7967
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 6380 7908 6776 7936
rect 4801 7871 4859 7877
rect 4801 7837 4813 7871
rect 4847 7837 4859 7871
rect 4801 7831 4859 7837
rect 5074 7828 5080 7880
rect 5132 7828 5138 7880
rect 5184 7868 5212 7896
rect 5353 7871 5411 7877
rect 5353 7868 5365 7871
rect 5184 7840 5365 7868
rect 5353 7837 5365 7840
rect 5399 7837 5411 7871
rect 5353 7831 5411 7837
rect 5626 7828 5632 7880
rect 5684 7868 5690 7880
rect 5902 7868 5908 7880
rect 5684 7840 5908 7868
rect 5684 7828 5690 7840
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6454 7868 6460 7880
rect 6288 7840 6460 7868
rect 5261 7803 5319 7809
rect 5261 7769 5273 7803
rect 5307 7800 5319 7803
rect 6288 7800 6316 7840
rect 6454 7828 6460 7840
rect 6512 7868 6518 7880
rect 6748 7877 6776 7908
rect 6840 7908 7665 7936
rect 6840 7877 6868 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 6641 7871 6699 7877
rect 6641 7868 6653 7871
rect 6512 7840 6653 7868
rect 6512 7828 6518 7840
rect 6641 7837 6653 7840
rect 6687 7837 6699 7871
rect 6641 7831 6699 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 5307 7772 6316 7800
rect 6365 7803 6423 7809
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 6365 7769 6377 7803
rect 6411 7769 6423 7803
rect 6656 7800 6684 7831
rect 7006 7828 7012 7880
rect 7064 7828 7070 7880
rect 7285 7803 7343 7809
rect 7285 7800 7297 7803
rect 6656 7772 7297 7800
rect 6365 7763 6423 7769
rect 7285 7769 7297 7772
rect 7331 7769 7343 7803
rect 7285 7763 7343 7769
rect 7469 7803 7527 7809
rect 7469 7769 7481 7803
rect 7515 7769 7527 7803
rect 7469 7763 7527 7769
rect 2501 7735 2559 7741
rect 2501 7701 2513 7735
rect 2547 7732 2559 7735
rect 4893 7735 4951 7741
rect 4893 7732 4905 7735
rect 2547 7704 4905 7732
rect 2547 7701 2559 7704
rect 2501 7695 2559 7701
rect 4893 7701 4905 7704
rect 4939 7732 4951 7735
rect 5350 7732 5356 7744
rect 4939 7704 5356 7732
rect 4939 7701 4951 7704
rect 4893 7695 4951 7701
rect 5350 7692 5356 7704
rect 5408 7732 5414 7744
rect 5445 7735 5503 7741
rect 5445 7732 5457 7735
rect 5408 7704 5457 7732
rect 5408 7692 5414 7704
rect 5445 7701 5457 7704
rect 5491 7701 5503 7735
rect 5445 7695 5503 7701
rect 5810 7692 5816 7744
rect 5868 7692 5874 7744
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6380 7732 6408 7763
rect 5960 7704 6408 7732
rect 6549 7735 6607 7741
rect 5960 7692 5966 7704
rect 6549 7701 6561 7735
rect 6595 7732 6607 7735
rect 7098 7732 7104 7744
rect 6595 7704 7104 7732
rect 6595 7701 6607 7704
rect 6549 7695 6607 7701
rect 7098 7692 7104 7704
rect 7156 7732 7162 7744
rect 7484 7732 7512 7763
rect 7156 7704 7512 7732
rect 7156 7692 7162 7704
rect 1104 7642 9108 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 4610 7642
rect 4662 7590 4674 7642
rect 4726 7590 4738 7642
rect 4790 7590 4802 7642
rect 4854 7590 4866 7642
rect 4918 7590 6610 7642
rect 6662 7590 6674 7642
rect 6726 7590 6738 7642
rect 6790 7590 6802 7642
rect 6854 7590 6866 7642
rect 6918 7590 8610 7642
rect 8662 7590 8674 7642
rect 8726 7590 8738 7642
rect 8790 7590 8802 7642
rect 8854 7590 8866 7642
rect 8918 7590 9108 7642
rect 1104 7568 9108 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 5074 7528 5080 7540
rect 3099 7500 5080 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 6454 7488 6460 7540
rect 6512 7488 6518 7540
rect 1854 7420 1860 7472
rect 1912 7460 1918 7472
rect 2498 7460 2504 7472
rect 1912 7432 2504 7460
rect 1912 7420 1918 7432
rect 2498 7420 2504 7432
rect 2556 7460 2562 7472
rect 2593 7463 2651 7469
rect 2593 7460 2605 7463
rect 2556 7432 2605 7460
rect 2556 7420 2562 7432
rect 2593 7429 2605 7432
rect 2639 7429 2651 7463
rect 5828 7460 5856 7488
rect 2593 7423 2651 7429
rect 4816 7432 5856 7460
rect 6472 7460 6500 7488
rect 6733 7463 6791 7469
rect 6472 7432 6684 7460
rect 4816 7401 4844 7432
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 5077 7395 5135 7401
rect 5077 7361 5089 7395
rect 5123 7392 5135 7395
rect 5166 7392 5172 7404
rect 5123 7364 5172 7392
rect 5123 7361 5135 7364
rect 5077 7355 5135 7361
rect 5166 7352 5172 7364
rect 5224 7352 5230 7404
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 5350 7392 5356 7404
rect 5307 7364 5356 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6656 7392 6684 7432
rect 6733 7429 6745 7463
rect 6779 7460 6791 7463
rect 6779 7432 7144 7460
rect 6779 7429 6791 7432
rect 6733 7423 6791 7429
rect 7116 7404 7144 7432
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6656 7364 6837 7392
rect 6549 7355 6607 7361
rect 6825 7361 6837 7364
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 6564 7324 6592 7355
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7392 8815 7395
rect 8803 7364 9260 7392
rect 8803 7361 8815 7364
rect 8757 7355 8815 7361
rect 9232 7336 9260 7364
rect 7282 7324 7288 7336
rect 6564 7296 7288 7324
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 1670 7216 1676 7268
rect 1728 7256 1734 7268
rect 2869 7259 2927 7265
rect 2869 7256 2881 7259
rect 1728 7228 2881 7256
rect 1728 7216 1734 7228
rect 2869 7225 2881 7228
rect 2915 7256 2927 7259
rect 2958 7256 2964 7268
rect 2915 7228 2964 7256
rect 2915 7225 2927 7228
rect 2869 7219 2927 7225
rect 2958 7216 2964 7228
rect 3016 7216 3022 7268
rect 4982 7216 4988 7268
rect 5040 7256 5046 7268
rect 8573 7259 8631 7265
rect 8573 7256 8585 7259
rect 5040 7228 8585 7256
rect 5040 7216 5046 7228
rect 8573 7225 8585 7228
rect 8619 7225 8631 7259
rect 8573 7219 8631 7225
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4580 7160 4629 7188
rect 4580 7148 4586 7160
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 4617 7151 4675 7157
rect 6365 7191 6423 7197
rect 6365 7157 6377 7191
rect 6411 7188 6423 7191
rect 6454 7188 6460 7200
rect 6411 7160 6460 7188
rect 6411 7157 6423 7160
rect 6365 7151 6423 7157
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 1104 7098 9108 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 3950 7098
rect 4002 7046 4014 7098
rect 4066 7046 4078 7098
rect 4130 7046 4142 7098
rect 4194 7046 4206 7098
rect 4258 7046 5950 7098
rect 6002 7046 6014 7098
rect 6066 7046 6078 7098
rect 6130 7046 6142 7098
rect 6194 7046 6206 7098
rect 6258 7046 7950 7098
rect 8002 7046 8014 7098
rect 8066 7046 8078 7098
rect 8130 7046 8142 7098
rect 8194 7046 8206 7098
rect 8258 7046 9108 7098
rect 1104 7024 9108 7046
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 7929 6987 7987 6993
rect 7929 6984 7941 6987
rect 7340 6956 7941 6984
rect 7340 6944 7346 6956
rect 7929 6953 7941 6956
rect 7975 6953 7987 6987
rect 7929 6947 7987 6953
rect 8021 6919 8079 6925
rect 8021 6885 8033 6919
rect 8067 6885 8079 6919
rect 8021 6879 8079 6885
rect 7834 6808 7840 6860
rect 7892 6848 7898 6860
rect 8036 6848 8064 6879
rect 7892 6820 8064 6848
rect 7892 6808 7898 6820
rect 8389 6715 8447 6721
rect 8389 6681 8401 6715
rect 8435 6712 8447 6715
rect 8478 6712 8484 6724
rect 8435 6684 8484 6712
rect 8435 6681 8447 6684
rect 8389 6675 8447 6681
rect 8478 6672 8484 6684
rect 8536 6672 8542 6724
rect 4154 6604 4160 6656
rect 4212 6644 4218 6656
rect 5350 6644 5356 6656
rect 4212 6616 5356 6644
rect 4212 6604 4218 6616
rect 5350 6604 5356 6616
rect 5408 6604 5414 6656
rect 1104 6554 9108 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 4610 6554
rect 4662 6502 4674 6554
rect 4726 6502 4738 6554
rect 4790 6502 4802 6554
rect 4854 6502 4866 6554
rect 4918 6502 6610 6554
rect 6662 6502 6674 6554
rect 6726 6502 6738 6554
rect 6790 6502 6802 6554
rect 6854 6502 6866 6554
rect 6918 6502 8610 6554
rect 8662 6502 8674 6554
rect 8726 6502 8738 6554
rect 8790 6502 8802 6554
rect 8854 6502 8866 6554
rect 8918 6502 9108 6554
rect 1104 6480 9108 6502
rect 1765 6443 1823 6449
rect 1765 6440 1777 6443
rect 1596 6412 1777 6440
rect 1596 6316 1624 6412
rect 1765 6409 1777 6412
rect 1811 6440 1823 6443
rect 2498 6440 2504 6452
rect 1811 6412 2504 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 2498 6400 2504 6412
rect 2556 6440 2562 6452
rect 2777 6443 2835 6449
rect 2556 6412 2636 6440
rect 2556 6400 2562 6412
rect 2608 6372 2636 6412
rect 2777 6409 2789 6443
rect 2823 6440 2835 6443
rect 2823 6412 4752 6440
rect 2823 6409 2835 6412
rect 2777 6403 2835 6409
rect 1688 6344 2452 6372
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 1688 6313 1716 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1820 6276 1961 6304
rect 1820 6264 1826 6276
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2041 6307 2099 6313
rect 2041 6273 2053 6307
rect 2087 6273 2099 6307
rect 2041 6267 2099 6273
rect 2056 6236 2084 6267
rect 2222 6264 2228 6316
rect 2280 6313 2286 6316
rect 2280 6304 2287 6313
rect 2280 6276 2325 6304
rect 2280 6267 2287 6276
rect 2280 6264 2286 6267
rect 2424 6245 2452 6344
rect 2608 6344 3096 6372
rect 2608 6313 2636 6344
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6273 2651 6307
rect 2869 6307 2927 6313
rect 2869 6304 2881 6307
rect 2593 6267 2651 6273
rect 2746 6276 2881 6304
rect 1780 6208 2084 6236
rect 2317 6239 2375 6245
rect 1780 6180 1808 6208
rect 2317 6205 2329 6239
rect 2363 6205 2375 6239
rect 2317 6199 2375 6205
rect 2409 6239 2467 6245
rect 2409 6205 2421 6239
rect 2455 6236 2467 6239
rect 2746 6236 2774 6276
rect 2869 6273 2881 6276
rect 2915 6304 2927 6307
rect 2958 6304 2964 6316
rect 2915 6276 2964 6304
rect 2915 6273 2927 6276
rect 2869 6267 2927 6273
rect 2958 6264 2964 6276
rect 3016 6264 3022 6316
rect 3068 6313 3096 6344
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3605 6307 3663 6313
rect 3605 6273 3617 6307
rect 3651 6304 3663 6307
rect 4154 6304 4160 6316
rect 3651 6276 4160 6304
rect 3651 6273 3663 6276
rect 3605 6267 3663 6273
rect 4154 6264 4160 6276
rect 4212 6264 4218 6316
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 4341 6307 4399 6313
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 4430 6304 4436 6316
rect 4387 6276 4436 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 2455 6208 2774 6236
rect 2455 6205 2467 6208
rect 2409 6199 2467 6205
rect 1762 6128 1768 6180
rect 1820 6128 1826 6180
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 1949 6171 2007 6177
rect 1949 6168 1961 6171
rect 1912 6140 1961 6168
rect 1912 6128 1918 6140
rect 1949 6137 1961 6140
rect 1995 6168 2007 6171
rect 2332 6168 2360 6199
rect 3694 6196 3700 6248
rect 3752 6236 3758 6248
rect 3878 6236 3884 6248
rect 3752 6208 3884 6236
rect 3752 6196 3758 6208
rect 3878 6196 3884 6208
rect 3936 6196 3942 6248
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4264 6236 4292 6267
rect 4430 6264 4436 6276
rect 4488 6264 4494 6316
rect 4522 6264 4528 6316
rect 4580 6264 4586 6316
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6304 4675 6307
rect 4724 6304 4752 6412
rect 5350 6400 5356 6452
rect 5408 6400 5414 6452
rect 7377 6443 7435 6449
rect 7377 6409 7389 6443
rect 7423 6409 7435 6443
rect 7377 6403 7435 6409
rect 4663 6276 4752 6304
rect 4985 6307 5043 6313
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5368 6304 5396 6400
rect 7098 6372 7104 6384
rect 6104 6344 7104 6372
rect 6104 6313 6132 6344
rect 7098 6332 7104 6344
rect 7156 6372 7162 6384
rect 7392 6372 7420 6403
rect 7156 6344 7420 6372
rect 7156 6332 7162 6344
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 8297 6375 8355 6381
rect 8297 6372 8309 6375
rect 7892 6344 8309 6372
rect 7892 6332 7898 6344
rect 8297 6341 8309 6344
rect 8343 6341 8355 6375
rect 8297 6335 8355 6341
rect 5031 6276 5396 6304
rect 6089 6307 6147 6313
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 6089 6273 6101 6307
rect 6135 6273 6147 6307
rect 6089 6267 6147 6273
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6304 7435 6307
rect 7466 6304 7472 6316
rect 7423 6276 7472 6304
rect 7423 6273 7435 6276
rect 7377 6267 7435 6273
rect 4019 6208 4292 6236
rect 4709 6239 4767 6245
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4709 6205 4721 6239
rect 4755 6205 4767 6239
rect 6380 6236 6408 6267
rect 4709 6199 4767 6205
rect 5828 6208 6408 6236
rect 6564 6236 6592 6267
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6304 8171 6307
rect 8478 6304 8484 6316
rect 8159 6276 8484 6304
rect 8159 6273 8171 6276
rect 8113 6267 8171 6273
rect 7576 6236 7604 6267
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 6564 6208 7941 6236
rect 1995 6140 2360 6168
rect 2961 6171 3019 6177
rect 1995 6137 2007 6140
rect 1949 6131 2007 6137
rect 2961 6137 2973 6171
rect 3007 6168 3019 6171
rect 4724 6168 4752 6199
rect 3007 6140 4752 6168
rect 4801 6171 4859 6177
rect 3007 6137 3019 6140
rect 2961 6131 3019 6137
rect 4801 6137 4813 6171
rect 4847 6168 4859 6171
rect 5828 6168 5856 6208
rect 6564 6168 6592 6208
rect 7929 6205 7941 6208
rect 7975 6205 7987 6239
rect 7929 6199 7987 6205
rect 4847 6140 5856 6168
rect 4847 6137 4859 6140
rect 4801 6131 4859 6137
rect 3418 6060 3424 6112
rect 3476 6100 3482 6112
rect 4065 6103 4123 6109
rect 4065 6100 4077 6103
rect 3476 6072 4077 6100
rect 3476 6060 3482 6072
rect 4065 6069 4077 6072
rect 4111 6069 4123 6103
rect 4065 6063 4123 6069
rect 4154 6060 4160 6112
rect 4212 6100 4218 6112
rect 4893 6103 4951 6109
rect 4893 6100 4905 6103
rect 4212 6072 4905 6100
rect 4212 6060 4218 6072
rect 4893 6069 4905 6072
rect 4939 6069 4951 6103
rect 4893 6063 4951 6069
rect 5442 6060 5448 6112
rect 5500 6100 5506 6112
rect 5828 6109 5856 6140
rect 6288 6140 6592 6168
rect 6288 6112 6316 6140
rect 5629 6103 5687 6109
rect 5629 6100 5641 6103
rect 5500 6072 5641 6100
rect 5500 6060 5506 6072
rect 5629 6069 5641 6072
rect 5675 6069 5687 6103
rect 5629 6063 5687 6069
rect 5813 6103 5871 6109
rect 5813 6069 5825 6103
rect 5859 6069 5871 6103
rect 5813 6063 5871 6069
rect 6270 6060 6276 6112
rect 6328 6060 6334 6112
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 6730 6100 6736 6112
rect 6503 6072 6736 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 6730 6060 6736 6072
rect 6788 6060 6794 6112
rect 1104 6010 9108 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 3950 6010
rect 4002 5958 4014 6010
rect 4066 5958 4078 6010
rect 4130 5958 4142 6010
rect 4194 5958 4206 6010
rect 4258 5958 5950 6010
rect 6002 5958 6014 6010
rect 6066 5958 6078 6010
rect 6130 5958 6142 6010
rect 6194 5958 6206 6010
rect 6258 5958 7950 6010
rect 8002 5958 8014 6010
rect 8066 5958 8078 6010
rect 8130 5958 8142 6010
rect 8194 5958 8206 6010
rect 8258 5958 9108 6010
rect 1104 5936 9108 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 1765 5899 1823 5905
rect 1765 5896 1777 5899
rect 1544 5868 1777 5896
rect 1544 5856 1550 5868
rect 1765 5865 1777 5868
rect 1811 5865 1823 5899
rect 1765 5859 1823 5865
rect 1854 5856 1860 5908
rect 1912 5856 1918 5908
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 7006 5896 7012 5908
rect 6779 5868 7012 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 7006 5856 7012 5868
rect 7064 5856 7070 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7116 5868 7941 5896
rect 1872 5760 1900 5856
rect 5166 5788 5172 5840
rect 5224 5828 5230 5840
rect 5224 5800 6592 5828
rect 5224 5788 5230 5800
rect 1949 5763 2007 5769
rect 1949 5760 1961 5763
rect 1872 5732 1961 5760
rect 1949 5729 1961 5732
rect 1995 5729 2007 5763
rect 5442 5760 5448 5772
rect 1949 5723 2007 5729
rect 5368 5732 5448 5760
rect 5368 5701 5396 5732
rect 5442 5720 5448 5732
rect 5500 5720 5506 5772
rect 5810 5760 5816 5772
rect 5736 5732 5816 5760
rect 5736 5701 5764 5732
rect 5810 5720 5816 5732
rect 5868 5760 5874 5772
rect 5868 5732 6500 5760
rect 5868 5720 5874 5732
rect 6270 5701 6276 5704
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5661 5411 5695
rect 5537 5695 5595 5701
rect 5537 5692 5549 5695
rect 5353 5655 5411 5661
rect 5460 5664 5549 5692
rect 1688 5624 1716 5655
rect 1854 5624 1860 5636
rect 1688 5596 1860 5624
rect 1854 5584 1860 5596
rect 1912 5584 1918 5636
rect 4430 5584 4436 5636
rect 4488 5624 4494 5636
rect 5460 5624 5488 5664
rect 5537 5661 5549 5664
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5629 5695 5687 5701
rect 5629 5661 5641 5695
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 5721 5695 5779 5701
rect 5721 5661 5733 5695
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5661 6147 5695
rect 6089 5655 6147 5661
rect 6237 5695 6276 5701
rect 6237 5661 6249 5695
rect 6237 5655 6276 5661
rect 4488 5596 5488 5624
rect 4488 5584 4494 5596
rect 5460 5568 5488 5596
rect 1762 5516 1768 5568
rect 1820 5556 1826 5568
rect 1949 5559 2007 5565
rect 1949 5556 1961 5559
rect 1820 5528 1961 5556
rect 1820 5516 1826 5528
rect 1949 5525 1961 5528
rect 1995 5525 2007 5559
rect 1949 5519 2007 5525
rect 5442 5516 5448 5568
rect 5500 5516 5506 5568
rect 5644 5556 5672 5655
rect 5997 5627 6055 5633
rect 5997 5593 6009 5627
rect 6043 5624 6055 5627
rect 6104 5624 6132 5655
rect 6270 5652 6276 5655
rect 6328 5652 6334 5704
rect 6472 5701 6500 5732
rect 6564 5701 6592 5800
rect 7116 5760 7144 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 7929 5859 7987 5865
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 8481 5831 8539 5837
rect 8481 5828 8493 5831
rect 7524 5800 8493 5828
rect 7524 5788 7530 5800
rect 7760 5769 7788 5800
rect 8481 5797 8493 5800
rect 8527 5797 8539 5831
rect 8481 5791 8539 5797
rect 6656 5732 7144 5760
rect 7745 5763 7803 5769
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5661 6515 5695
rect 6457 5655 6515 5661
rect 6554 5695 6612 5701
rect 6554 5661 6566 5695
rect 6600 5661 6612 5695
rect 6554 5655 6612 5661
rect 6043 5596 6132 5624
rect 6043 5593 6055 5596
rect 5997 5587 6055 5593
rect 6362 5584 6368 5636
rect 6420 5584 6426 5636
rect 6472 5624 6500 5655
rect 6656 5624 6684 5732
rect 7745 5729 7757 5763
rect 7791 5729 7803 5763
rect 7745 5723 7803 5729
rect 8128 5732 8432 5760
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 6788 5664 7573 5692
rect 6788 5652 6794 5664
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 8128 5701 8156 5732
rect 8404 5701 8432 5732
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 7892 5664 8125 5692
rect 7892 5652 7898 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8297 5695 8355 5701
rect 8297 5661 8309 5695
rect 8343 5661 8355 5695
rect 8297 5655 8355 5661
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 6472 5596 6684 5624
rect 6748 5556 6776 5652
rect 8312 5624 8340 5655
rect 8478 5652 8484 5704
rect 8536 5692 8542 5704
rect 8573 5695 8631 5701
rect 8573 5692 8585 5695
rect 8536 5664 8585 5692
rect 8536 5652 8542 5664
rect 8573 5661 8585 5664
rect 8619 5661 8631 5695
rect 8573 5655 8631 5661
rect 8496 5624 8524 5652
rect 8312 5596 8524 5624
rect 5644 5528 6776 5556
rect 7374 5516 7380 5568
rect 7432 5516 7438 5568
rect 1104 5466 9108 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 4610 5466
rect 4662 5414 4674 5466
rect 4726 5414 4738 5466
rect 4790 5414 4802 5466
rect 4854 5414 4866 5466
rect 4918 5414 6610 5466
rect 6662 5414 6674 5466
rect 6726 5414 6738 5466
rect 6790 5414 6802 5466
rect 6854 5414 6866 5466
rect 6918 5414 8610 5466
rect 8662 5414 8674 5466
rect 8726 5414 8738 5466
rect 8790 5414 8802 5466
rect 8854 5414 8866 5466
rect 8918 5414 9108 5466
rect 1104 5392 9108 5414
rect 2774 5312 2780 5364
rect 2832 5352 2838 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 2832 5324 3157 5352
rect 2832 5312 2838 5324
rect 3145 5321 3157 5324
rect 3191 5352 3203 5355
rect 3326 5352 3332 5364
rect 3191 5324 3332 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3326 5312 3332 5324
rect 3384 5352 3390 5364
rect 3786 5352 3792 5364
rect 3384 5324 3792 5352
rect 3384 5312 3390 5324
rect 3786 5312 3792 5324
rect 3844 5312 3850 5364
rect 4985 5355 5043 5361
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 6362 5352 6368 5364
rect 5031 5324 6368 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 934 5244 940 5296
rect 992 5284 998 5296
rect 1397 5287 1455 5293
rect 1397 5284 1409 5287
rect 992 5256 1409 5284
rect 992 5244 998 5256
rect 1397 5253 1409 5256
rect 1443 5253 1455 5287
rect 1397 5247 1455 5253
rect 1765 5287 1823 5293
rect 1765 5253 1777 5287
rect 1811 5284 1823 5287
rect 3418 5284 3424 5296
rect 1811 5256 3424 5284
rect 1811 5253 1823 5256
rect 1765 5247 1823 5253
rect 3418 5244 3424 5256
rect 3476 5244 3482 5296
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5216 3295 5219
rect 3602 5216 3608 5228
rect 3283 5188 3608 5216
rect 3283 5185 3295 5188
rect 3237 5179 3295 5185
rect 3252 5092 3280 5179
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 5074 5176 5080 5228
rect 5132 5176 5138 5228
rect 5261 5219 5319 5225
rect 5261 5185 5273 5219
rect 5307 5216 5319 5219
rect 5810 5216 5816 5228
rect 5307 5188 5816 5216
rect 5307 5185 5319 5188
rect 5261 5179 5319 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 3234 5040 3240 5092
rect 3292 5040 3298 5092
rect 4798 4972 4804 5024
rect 4856 4972 4862 5024
rect 1104 4922 9108 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 3950 4922
rect 4002 4870 4014 4922
rect 4066 4870 4078 4922
rect 4130 4870 4142 4922
rect 4194 4870 4206 4922
rect 4258 4870 5950 4922
rect 6002 4870 6014 4922
rect 6066 4870 6078 4922
rect 6130 4870 6142 4922
rect 6194 4870 6206 4922
rect 6258 4870 7950 4922
rect 8002 4870 8014 4922
rect 8066 4870 8078 4922
rect 8130 4870 8142 4922
rect 8194 4870 8206 4922
rect 8258 4870 9108 4922
rect 1104 4848 9108 4870
rect 1486 4768 1492 4820
rect 1544 4768 1550 4820
rect 1670 4768 1676 4820
rect 1728 4808 1734 4820
rect 2317 4811 2375 4817
rect 2317 4808 2329 4811
rect 1728 4780 2329 4808
rect 1728 4768 1734 4780
rect 2317 4777 2329 4780
rect 2363 4808 2375 4811
rect 2406 4808 2412 4820
rect 2363 4780 2412 4808
rect 2363 4777 2375 4780
rect 2317 4771 2375 4777
rect 2406 4768 2412 4780
rect 2464 4768 2470 4820
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2516 4780 2973 4808
rect 1504 4672 1532 4768
rect 2516 4681 2544 4780
rect 2961 4777 2973 4780
rect 3007 4808 3019 4811
rect 3418 4808 3424 4820
rect 3007 4780 3424 4808
rect 3007 4777 3019 4780
rect 2961 4771 3019 4777
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3651 4780 3985 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3973 4777 3985 4780
rect 4019 4808 4031 4811
rect 4019 4780 4384 4808
rect 4019 4777 4031 4780
rect 3973 4771 4031 4777
rect 3145 4743 3203 4749
rect 3145 4709 3157 4743
rect 3191 4709 3203 4743
rect 3145 4703 3203 4709
rect 2501 4675 2559 4681
rect 2501 4672 2513 4675
rect 1504 4644 2513 4672
rect 1854 4564 1860 4616
rect 1912 4564 1918 4616
rect 1964 4613 1992 4644
rect 2501 4641 2513 4644
rect 2547 4641 2559 4675
rect 3160 4672 3188 4703
rect 4356 4681 4384 4780
rect 5074 4768 5080 4820
rect 5132 4768 5138 4820
rect 4522 4700 4528 4752
rect 4580 4740 4586 4752
rect 4617 4743 4675 4749
rect 4617 4740 4629 4743
rect 4580 4712 4629 4740
rect 4580 4700 4586 4712
rect 4617 4709 4629 4712
rect 4663 4709 4675 4743
rect 4617 4703 4675 4709
rect 4801 4743 4859 4749
rect 4801 4709 4813 4743
rect 4847 4740 4859 4743
rect 4890 4740 4896 4752
rect 4847 4712 4896 4740
rect 4847 4709 4859 4712
rect 4801 4703 4859 4709
rect 4890 4700 4896 4712
rect 4948 4700 4954 4752
rect 4341 4675 4399 4681
rect 3160 4644 4292 4672
rect 2501 4635 2559 4641
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4573 2007 4607
rect 1949 4567 2007 4573
rect 2225 4607 2283 4613
rect 2225 4573 2237 4607
rect 2271 4573 2283 4607
rect 2225 4567 2283 4573
rect 1872 4536 1900 4564
rect 2240 4536 2268 4567
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 2884 4604 3020 4606
rect 3050 4604 3056 4616
rect 2464 4578 3056 4604
rect 2464 4576 2912 4578
rect 2464 4564 2470 4576
rect 2992 4573 3056 4578
rect 2774 4536 2780 4548
rect 1872 4508 2780 4536
rect 2774 4496 2780 4508
rect 2832 4536 2838 4548
rect 2992 4542 3019 4573
rect 3007 4539 3019 4542
rect 3053 4564 3056 4573
rect 3108 4604 3114 4616
rect 3237 4607 3295 4613
rect 3237 4604 3249 4607
rect 3108 4576 3249 4604
rect 3108 4564 3114 4576
rect 3237 4573 3249 4576
rect 3283 4573 3295 4607
rect 3237 4567 3295 4573
rect 3326 4564 3332 4616
rect 3384 4564 3390 4616
rect 4264 4604 4292 4644
rect 4341 4641 4353 4675
rect 4387 4672 4399 4675
rect 5092 4672 5120 4768
rect 4387 4644 5120 4672
rect 4387 4641 4399 4644
rect 4341 4635 4399 4641
rect 4798 4604 4804 4616
rect 4264 4576 4804 4604
rect 4798 4564 4804 4576
rect 4856 4604 4862 4616
rect 5077 4607 5135 4613
rect 5077 4604 5089 4607
rect 4856 4576 5089 4604
rect 4856 4564 4862 4576
rect 5077 4573 5089 4576
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5626 4564 5632 4616
rect 5684 4604 5690 4616
rect 5902 4604 5908 4616
rect 5684 4576 5908 4604
rect 5684 4564 5690 4576
rect 5902 4564 5908 4576
rect 5960 4564 5966 4616
rect 3053 4542 3091 4564
rect 3053 4539 3065 4542
rect 2832 4508 2877 4536
rect 3007 4533 3065 4539
rect 2832 4496 2838 4508
rect 3786 4496 3792 4548
rect 3844 4536 3850 4548
rect 3844 4508 4752 4536
rect 3844 4496 3850 4508
rect 2130 4428 2136 4480
rect 2188 4428 2194 4480
rect 2501 4471 2559 4477
rect 2501 4437 2513 4471
rect 2547 4468 2559 4471
rect 3989 4471 4047 4477
rect 3989 4468 4001 4471
rect 2547 4440 4001 4468
rect 2547 4437 2559 4440
rect 2501 4431 2559 4437
rect 3989 4437 4001 4440
rect 4035 4437 4047 4471
rect 3989 4431 4047 4437
rect 4154 4428 4160 4480
rect 4212 4428 4218 4480
rect 4724 4468 4752 4508
rect 4890 4496 4896 4548
rect 4948 4496 4954 4548
rect 5644 4536 5672 4564
rect 5000 4508 5672 4536
rect 5000 4468 5028 4508
rect 4724 4440 5028 4468
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4468 5319 4471
rect 6362 4468 6368 4480
rect 5307 4440 6368 4468
rect 5307 4437 5319 4440
rect 5261 4431 5319 4437
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 1104 4378 9108 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 4610 4378
rect 4662 4326 4674 4378
rect 4726 4326 4738 4378
rect 4790 4326 4802 4378
rect 4854 4326 4866 4378
rect 4918 4326 6610 4378
rect 6662 4326 6674 4378
rect 6726 4326 6738 4378
rect 6790 4326 6802 4378
rect 6854 4326 6866 4378
rect 6918 4326 8610 4378
rect 8662 4326 8674 4378
rect 8726 4326 8738 4378
rect 8790 4326 8802 4378
rect 8854 4326 8866 4378
rect 8918 4326 9108 4378
rect 1104 4304 9108 4326
rect 3237 4267 3295 4273
rect 3237 4233 3249 4267
rect 3283 4264 3295 4267
rect 3786 4264 3792 4276
rect 3283 4236 3792 4264
rect 3283 4233 3295 4236
rect 3237 4227 3295 4233
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 4154 4224 4160 4276
rect 4212 4264 4218 4276
rect 5442 4264 5448 4276
rect 4212 4236 5448 4264
rect 4212 4224 4218 4236
rect 5442 4224 5448 4236
rect 5500 4264 5506 4276
rect 5500 4236 6684 4264
rect 5500 4224 5506 4236
rect 2130 4156 2136 4208
rect 2188 4196 2194 4208
rect 5166 4196 5172 4208
rect 2188 4168 5172 4196
rect 2188 4156 2194 4168
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 5902 4156 5908 4208
rect 5960 4156 5966 4208
rect 6365 4199 6423 4205
rect 6365 4165 6377 4199
rect 6411 4196 6423 4199
rect 6454 4196 6460 4208
rect 6411 4168 6460 4196
rect 6411 4165 6423 4168
rect 6365 4159 6423 4165
rect 3050 4088 3056 4140
rect 3108 4088 3114 4140
rect 5327 4131 5385 4137
rect 5327 4097 5339 4131
rect 5373 4097 5385 4131
rect 5327 4091 5385 4097
rect 3234 4020 3240 4072
rect 3292 4060 3298 4072
rect 3421 4063 3479 4069
rect 3421 4060 3433 4063
rect 3292 4032 3433 4060
rect 3292 4020 3298 4032
rect 3421 4029 3433 4032
rect 3467 4060 3479 4063
rect 4890 4060 4896 4072
rect 3467 4032 4896 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 4890 4020 4896 4032
rect 4948 4020 4954 4072
rect 5074 4020 5080 4072
rect 5132 4060 5138 4072
rect 5169 4063 5227 4069
rect 5169 4060 5181 4063
rect 5132 4032 5181 4060
rect 5132 4020 5138 4032
rect 5169 4029 5181 4032
rect 5215 4029 5227 4063
rect 5169 4023 5227 4029
rect 3418 3884 3424 3936
rect 3476 3884 3482 3936
rect 5342 3924 5370 4091
rect 5442 4088 5448 4140
rect 5500 4088 5506 4140
rect 5537 4131 5595 4137
rect 5537 4097 5549 4131
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5629 4131 5687 4137
rect 5629 4097 5641 4131
rect 5675 4097 5687 4131
rect 5629 4091 5687 4097
rect 6089 4131 6147 4137
rect 6089 4097 6101 4131
rect 6135 4097 6147 4131
rect 6089 4091 6147 4097
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4128 6239 4131
rect 6380 4128 6408 4159
rect 6454 4156 6460 4168
rect 6512 4156 6518 4208
rect 6227 4100 6408 4128
rect 6549 4131 6607 4137
rect 6227 4097 6239 4100
rect 6181 4091 6239 4097
rect 6549 4097 6561 4131
rect 6595 4097 6607 4131
rect 6656 4128 6684 4236
rect 7484 4168 7696 4196
rect 7193 4131 7251 4137
rect 7193 4128 7205 4131
rect 6656 4100 7205 4128
rect 6549 4091 6607 4097
rect 7193 4097 7205 4100
rect 7239 4097 7251 4131
rect 7193 4091 7251 4097
rect 5552 4004 5580 4091
rect 5644 4060 5672 4091
rect 6104 4060 6132 4091
rect 6270 4060 6276 4072
rect 5644 4032 6040 4060
rect 6104 4032 6276 4060
rect 5534 3952 5540 4004
rect 5592 3952 5598 4004
rect 5905 3995 5963 4001
rect 5905 3992 5917 3995
rect 5737 3964 5917 3992
rect 5737 3936 5765 3964
rect 5905 3961 5917 3964
rect 5951 3961 5963 3995
rect 6012 3992 6040 4032
rect 6270 4020 6276 4032
rect 6328 4060 6334 4072
rect 6564 4060 6592 4091
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7484 4128 7512 4168
rect 7432 4100 7512 4128
rect 7432 4088 7438 4100
rect 7558 4088 7564 4140
rect 7616 4088 7622 4140
rect 7668 4128 7696 4168
rect 7745 4131 7803 4137
rect 7745 4128 7757 4131
rect 7668 4100 7757 4128
rect 7745 4097 7757 4100
rect 7791 4097 7803 4131
rect 7745 4091 7803 4097
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 6328 4032 7481 4060
rect 6328 4020 6334 4032
rect 7469 4029 7481 4032
rect 7515 4029 7527 4063
rect 7469 4023 7527 4029
rect 7653 3995 7711 4001
rect 7653 3992 7665 3995
rect 6012 3964 7665 3992
rect 5905 3955 5963 3961
rect 7653 3961 7665 3964
rect 7699 3961 7711 3995
rect 7653 3955 7711 3961
rect 5718 3924 5724 3936
rect 5342 3896 5724 3924
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 5813 3927 5871 3933
rect 5813 3893 5825 3927
rect 5859 3924 5871 3927
rect 5994 3924 6000 3936
rect 5859 3896 6000 3924
rect 5859 3893 5871 3896
rect 5813 3887 5871 3893
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6730 3884 6736 3936
rect 6788 3884 6794 3936
rect 7006 3884 7012 3936
rect 7064 3884 7070 3936
rect 1104 3834 9108 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 3950 3834
rect 4002 3782 4014 3834
rect 4066 3782 4078 3834
rect 4130 3782 4142 3834
rect 4194 3782 4206 3834
rect 4258 3782 5950 3834
rect 6002 3782 6014 3834
rect 6066 3782 6078 3834
rect 6130 3782 6142 3834
rect 6194 3782 6206 3834
rect 6258 3782 7950 3834
rect 8002 3782 8014 3834
rect 8066 3782 8078 3834
rect 8130 3782 8142 3834
rect 8194 3782 8206 3834
rect 8258 3782 9108 3834
rect 1104 3760 9108 3782
rect 6086 3720 6092 3732
rect 5552 3692 6092 3720
rect 4522 3612 4528 3664
rect 4580 3652 4586 3664
rect 5552 3652 5580 3692
rect 6086 3680 6092 3692
rect 6144 3720 6150 3732
rect 7558 3720 7564 3732
rect 6144 3692 7564 3720
rect 6144 3680 6150 3692
rect 7558 3680 7564 3692
rect 7616 3680 7622 3732
rect 8573 3655 8631 3661
rect 8573 3652 8585 3655
rect 4580 3624 5580 3652
rect 5644 3624 8585 3652
rect 4580 3612 4586 3624
rect 4890 3544 4896 3596
rect 4948 3584 4954 3596
rect 5644 3584 5672 3624
rect 8573 3621 8585 3624
rect 8619 3621 8631 3655
rect 8573 3615 8631 3621
rect 6362 3584 6368 3596
rect 4948 3556 5672 3584
rect 5920 3556 6368 3584
rect 4948 3544 4954 3556
rect 5534 3476 5540 3528
rect 5592 3476 5598 3528
rect 5626 3476 5632 3528
rect 5684 3476 5690 3528
rect 5722 3519 5780 3525
rect 5722 3485 5734 3519
rect 5768 3485 5780 3519
rect 5722 3479 5780 3485
rect 5552 3448 5580 3476
rect 5736 3448 5764 3479
rect 5810 3448 5816 3460
rect 5552 3420 5816 3448
rect 5810 3408 5816 3420
rect 5868 3408 5874 3460
rect 5920 3457 5948 3556
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 6730 3544 6736 3596
rect 6788 3544 6794 3596
rect 6135 3519 6193 3525
rect 6135 3485 6147 3519
rect 6181 3516 6193 3519
rect 6748 3516 6776 3544
rect 6181 3488 6776 3516
rect 8757 3519 8815 3525
rect 6181 3485 6193 3488
rect 6135 3479 6193 3485
rect 8757 3485 8769 3519
rect 8803 3516 8815 3519
rect 9214 3516 9220 3528
rect 8803 3488 9220 3516
rect 8803 3485 8815 3488
rect 8757 3479 8815 3485
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 5905 3451 5963 3457
rect 5905 3417 5917 3451
rect 5951 3417 5963 3451
rect 5905 3411 5963 3417
rect 5997 3451 6055 3457
rect 5997 3417 6009 3451
rect 6043 3417 6055 3451
rect 5997 3411 6055 3417
rect 5718 3340 5724 3392
rect 5776 3380 5782 3392
rect 6012 3380 6040 3411
rect 5776 3352 6040 3380
rect 5776 3340 5782 3352
rect 6270 3340 6276 3392
rect 6328 3340 6334 3392
rect 1104 3290 9108 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 4610 3290
rect 4662 3238 4674 3290
rect 4726 3238 4738 3290
rect 4790 3238 4802 3290
rect 4854 3238 4866 3290
rect 4918 3238 6610 3290
rect 6662 3238 6674 3290
rect 6726 3238 6738 3290
rect 6790 3238 6802 3290
rect 6854 3238 6866 3290
rect 6918 3238 8610 3290
rect 8662 3238 8674 3290
rect 8726 3238 8738 3290
rect 8790 3238 8802 3290
rect 8854 3238 8866 3290
rect 8918 3238 9108 3290
rect 1104 3216 9108 3238
rect 4157 3179 4215 3185
rect 4157 3145 4169 3179
rect 4203 3176 4215 3179
rect 4522 3176 4528 3188
rect 4203 3148 4528 3176
rect 4203 3145 4215 3148
rect 4157 3139 4215 3145
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 4893 3179 4951 3185
rect 4893 3145 4905 3179
rect 4939 3176 4951 3179
rect 5074 3176 5080 3188
rect 4939 3148 5080 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5166 3136 5172 3188
rect 5224 3185 5230 3188
rect 5224 3179 5243 3185
rect 5231 3145 5243 3179
rect 5224 3139 5243 3145
rect 5353 3179 5411 3185
rect 5353 3145 5365 3179
rect 5399 3176 5411 3179
rect 5626 3176 5632 3188
rect 5399 3148 5632 3176
rect 5399 3145 5411 3148
rect 5353 3139 5411 3145
rect 5224 3136 5230 3139
rect 5626 3136 5632 3148
rect 5684 3136 5690 3188
rect 5810 3136 5816 3188
rect 5868 3136 5874 3188
rect 6086 3136 6092 3188
rect 6144 3136 6150 3188
rect 6178 3136 6184 3188
rect 6236 3136 6242 3188
rect 7374 3136 7380 3188
rect 7432 3136 7438 3188
rect 1765 3111 1823 3117
rect 1765 3077 1777 3111
rect 1811 3108 1823 3111
rect 3142 3108 3148 3120
rect 1811 3080 3148 3108
rect 1811 3077 1823 3080
rect 1765 3071 1823 3077
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 4985 3111 5043 3117
rect 4985 3108 4997 3111
rect 4172 3080 4997 3108
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 4172 3049 4200 3080
rect 4985 3077 4997 3080
rect 5031 3108 5043 3111
rect 5031 3080 5672 3108
rect 5031 3077 5043 3080
rect 4985 3071 5043 3077
rect 5644 3049 5672 3080
rect 4157 3043 4215 3049
rect 4157 3040 4169 3043
rect 2924 3012 4169 3040
rect 2924 3000 2930 3012
rect 4157 3009 4169 3012
rect 4203 3009 4215 3043
rect 4157 3003 4215 3009
rect 4341 3043 4399 3049
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4387 3012 4445 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 4433 3003 4491 3009
rect 5184 3012 5457 3040
rect 934 2796 940 2848
rect 992 2836 998 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 992 2808 1501 2836
rect 992 2796 998 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 4172 2836 4200 3003
rect 4448 2972 4476 3003
rect 5184 2972 5212 3012
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5629 3043 5687 3049
rect 5629 3009 5641 3043
rect 5675 3009 5687 3043
rect 5828 3040 5856 3136
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5828 3012 6009 3040
rect 5629 3003 5687 3009
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 6104 3040 6132 3136
rect 6196 3108 6224 3136
rect 6196 3080 7236 3108
rect 6181 3043 6239 3049
rect 6181 3040 6193 3043
rect 6104 3012 6193 3040
rect 5997 3003 6055 3009
rect 6181 3009 6193 3012
rect 6227 3009 6239 3043
rect 6181 3003 6239 3009
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 6328 3012 6653 3040
rect 6328 3000 6334 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 6641 3003 6699 3009
rect 6825 3043 6883 3049
rect 6825 3009 6837 3043
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3040 6975 3043
rect 7006 3040 7012 3052
rect 6963 3012 7012 3040
rect 6963 3009 6975 3012
rect 6917 3003 6975 3009
rect 4448 2944 5212 2972
rect 6840 2972 6868 3003
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7208 3049 7236 3080
rect 7392 3049 7420 3136
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 7377 3043 7435 3049
rect 7377 3009 7389 3043
rect 7423 3009 7435 3043
rect 7377 3003 7435 3009
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 6840 2944 7297 2972
rect 5184 2845 5212 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 7190 2904 7196 2916
rect 5828 2876 7196 2904
rect 4525 2839 4583 2845
rect 4525 2836 4537 2839
rect 4172 2808 4537 2836
rect 1489 2799 1547 2805
rect 4525 2805 4537 2808
rect 4571 2805 4583 2839
rect 4525 2799 4583 2805
rect 5169 2839 5227 2845
rect 5169 2805 5181 2839
rect 5215 2836 5227 2839
rect 5828 2836 5856 2876
rect 7190 2864 7196 2876
rect 7248 2864 7254 2916
rect 5215 2808 5856 2836
rect 5215 2805 5227 2808
rect 5169 2799 5227 2805
rect 6454 2796 6460 2848
rect 6512 2796 6518 2848
rect 1104 2746 9108 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 3950 2746
rect 4002 2694 4014 2746
rect 4066 2694 4078 2746
rect 4130 2694 4142 2746
rect 4194 2694 4206 2746
rect 4258 2694 5950 2746
rect 6002 2694 6014 2746
rect 6066 2694 6078 2746
rect 6130 2694 6142 2746
rect 6194 2694 6206 2746
rect 6258 2694 7950 2746
rect 8002 2694 8014 2746
rect 8066 2694 8078 2746
rect 8130 2694 8142 2746
rect 8194 2694 8206 2746
rect 8258 2694 9108 2746
rect 1104 2672 9108 2694
rect 1578 2592 1584 2644
rect 1636 2592 1642 2644
rect 2866 2592 2872 2644
rect 2924 2592 2930 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 7248 2604 8217 2632
rect 7248 2592 7254 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 8205 2595 8263 2601
rect 8478 2592 8484 2644
rect 8536 2632 8542 2644
rect 8665 2635 8723 2641
rect 8665 2632 8677 2635
rect 8536 2604 8677 2632
rect 8536 2592 8542 2604
rect 8665 2601 8677 2604
rect 8711 2601 8723 2635
rect 8665 2595 8723 2601
rect 2682 2388 2688 2440
rect 2740 2388 2746 2440
rect 5445 2431 5503 2437
rect 5445 2397 5457 2431
rect 5491 2428 5503 2431
rect 6454 2428 6460 2440
rect 5491 2400 6460 2428
rect 5491 2397 5503 2400
rect 5445 2391 5503 2397
rect 6454 2388 6460 2400
rect 6512 2388 6518 2440
rect 8389 2431 8447 2437
rect 8389 2397 8401 2431
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 72 2332 1501 2360
rect 72 2320 78 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 8404 2360 8432 2391
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 8404 2332 9076 2360
rect 1489 2323 1547 2329
rect 9048 2304 9076 2332
rect 5166 2252 5172 2304
rect 5224 2252 5230 2304
rect 9030 2252 9036 2304
rect 9088 2252 9094 2304
rect 1104 2202 9108 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 4610 2202
rect 4662 2150 4674 2202
rect 4726 2150 4738 2202
rect 4790 2150 4802 2202
rect 4854 2150 4866 2202
rect 4918 2150 6610 2202
rect 6662 2150 6674 2202
rect 6726 2150 6738 2202
rect 6790 2150 6802 2202
rect 6854 2150 6866 2202
rect 6918 2150 8610 2202
rect 8662 2150 8674 2202
rect 8726 2150 8738 2202
rect 8790 2150 8802 2202
rect 8854 2150 8866 2202
rect 8918 2150 9108 2202
rect 1104 2128 9108 2150
<< via1 >>
rect 2610 9766 2662 9818
rect 2674 9766 2726 9818
rect 2738 9766 2790 9818
rect 2802 9766 2854 9818
rect 2866 9766 2918 9818
rect 4610 9766 4662 9818
rect 4674 9766 4726 9818
rect 4738 9766 4790 9818
rect 4802 9766 4854 9818
rect 4866 9766 4918 9818
rect 6610 9766 6662 9818
rect 6674 9766 6726 9818
rect 6738 9766 6790 9818
rect 6802 9766 6854 9818
rect 6866 9766 6918 9818
rect 8610 9766 8662 9818
rect 8674 9766 8726 9818
rect 8738 9766 8790 9818
rect 8802 9766 8854 9818
rect 8866 9766 8918 9818
rect 1308 9596 1360 9648
rect 1860 9639 1912 9648
rect 1860 9605 1869 9639
rect 1869 9605 1903 9639
rect 1903 9605 1912 9639
rect 1860 9596 1912 9605
rect 4528 9596 4580 9648
rect 7380 9596 7432 9648
rect 7748 9596 7800 9648
rect 9680 9596 9732 9648
rect 7288 9571 7340 9580
rect 7288 9537 7297 9571
rect 7297 9537 7331 9571
rect 7331 9537 7340 9571
rect 7288 9528 7340 9537
rect 8944 9528 8996 9580
rect 1492 9324 1544 9376
rect 1676 9324 1728 9376
rect 4988 9324 5040 9376
rect 7840 9324 7892 9376
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 3950 9222 4002 9274
rect 4014 9222 4066 9274
rect 4078 9222 4130 9274
rect 4142 9222 4194 9274
rect 4206 9222 4258 9274
rect 5950 9222 6002 9274
rect 6014 9222 6066 9274
rect 6078 9222 6130 9274
rect 6142 9222 6194 9274
rect 6206 9222 6258 9274
rect 7950 9222 8002 9274
rect 8014 9222 8066 9274
rect 8078 9222 8130 9274
rect 8142 9222 8194 9274
rect 8206 9222 8258 9274
rect 7288 9120 7340 9172
rect 940 8916 992 8968
rect 1768 8916 1820 8968
rect 1492 8848 1544 8900
rect 3516 8984 3568 9036
rect 4160 8916 4212 8968
rect 5724 8916 5776 8968
rect 3332 8780 3384 8832
rect 3424 8780 3476 8832
rect 3608 8823 3660 8832
rect 3608 8789 3617 8823
rect 3617 8789 3651 8823
rect 3651 8789 3660 8823
rect 3608 8780 3660 8789
rect 3700 8780 3752 8832
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 4610 8678 4662 8730
rect 4674 8678 4726 8730
rect 4738 8678 4790 8730
rect 4802 8678 4854 8730
rect 4866 8678 4918 8730
rect 6610 8678 6662 8730
rect 6674 8678 6726 8730
rect 6738 8678 6790 8730
rect 6802 8678 6854 8730
rect 6866 8678 6918 8730
rect 8610 8678 8662 8730
rect 8674 8678 8726 8730
rect 8738 8678 8790 8730
rect 8802 8678 8854 8730
rect 8866 8678 8918 8730
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 3240 8576 3292 8628
rect 3608 8619 3660 8628
rect 3608 8585 3635 8619
rect 3635 8585 3660 8619
rect 3608 8576 3660 8585
rect 4988 8576 5040 8628
rect 3792 8551 3844 8560
rect 3792 8517 3801 8551
rect 3801 8517 3835 8551
rect 3835 8517 3844 8551
rect 3792 8508 3844 8517
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 3332 8483 3384 8492
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 4160 8483 4212 8492
rect 4160 8449 4169 8483
rect 4169 8449 4203 8483
rect 4203 8449 4212 8483
rect 4160 8440 4212 8449
rect 3148 8304 3200 8356
rect 3700 8304 3752 8356
rect 2964 8236 3016 8288
rect 3516 8236 3568 8288
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 5172 8279 5224 8288
rect 5172 8245 5181 8279
rect 5181 8245 5215 8279
rect 5215 8245 5224 8279
rect 5172 8236 5224 8245
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 3950 8134 4002 8186
rect 4014 8134 4066 8186
rect 4078 8134 4130 8186
rect 4142 8134 4194 8186
rect 4206 8134 4258 8186
rect 5950 8134 6002 8186
rect 6014 8134 6066 8186
rect 6078 8134 6130 8186
rect 6142 8134 6194 8186
rect 6206 8134 6258 8186
rect 7950 8134 8002 8186
rect 8014 8134 8066 8186
rect 8078 8134 8130 8186
rect 8142 8134 8194 8186
rect 8206 8134 8258 8186
rect 7748 8032 7800 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 1860 7871 1912 7880
rect 1860 7837 1869 7871
rect 1869 7837 1903 7871
rect 1903 7837 1912 7871
rect 1860 7828 1912 7837
rect 5172 7896 5224 7948
rect 5080 7871 5132 7880
rect 5080 7837 5089 7871
rect 5089 7837 5123 7871
rect 5123 7837 5132 7871
rect 5080 7828 5132 7837
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 5908 7828 5960 7880
rect 6460 7828 6512 7880
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 5356 7692 5408 7744
rect 5816 7735 5868 7744
rect 5816 7701 5825 7735
rect 5825 7701 5859 7735
rect 5859 7701 5868 7735
rect 5816 7692 5868 7701
rect 5908 7692 5960 7744
rect 7104 7692 7156 7744
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 4610 7590 4662 7642
rect 4674 7590 4726 7642
rect 4738 7590 4790 7642
rect 4802 7590 4854 7642
rect 4866 7590 4918 7642
rect 6610 7590 6662 7642
rect 6674 7590 6726 7642
rect 6738 7590 6790 7642
rect 6802 7590 6854 7642
rect 6866 7590 6918 7642
rect 8610 7590 8662 7642
rect 8674 7590 8726 7642
rect 8738 7590 8790 7642
rect 8802 7590 8854 7642
rect 8866 7590 8918 7642
rect 5080 7488 5132 7540
rect 5816 7488 5868 7540
rect 6460 7488 6512 7540
rect 1860 7420 1912 7472
rect 2504 7420 2556 7472
rect 5172 7352 5224 7404
rect 5356 7352 5408 7404
rect 7104 7352 7156 7404
rect 7288 7284 7340 7336
rect 9220 7284 9272 7336
rect 1676 7216 1728 7268
rect 2964 7216 3016 7268
rect 4988 7216 5040 7268
rect 4528 7148 4580 7200
rect 6460 7148 6512 7200
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 3950 7046 4002 7098
rect 4014 7046 4066 7098
rect 4078 7046 4130 7098
rect 4142 7046 4194 7098
rect 4206 7046 4258 7098
rect 5950 7046 6002 7098
rect 6014 7046 6066 7098
rect 6078 7046 6130 7098
rect 6142 7046 6194 7098
rect 6206 7046 6258 7098
rect 7950 7046 8002 7098
rect 8014 7046 8066 7098
rect 8078 7046 8130 7098
rect 8142 7046 8194 7098
rect 8206 7046 8258 7098
rect 7288 6944 7340 6996
rect 7840 6808 7892 6860
rect 8484 6672 8536 6724
rect 4160 6604 4212 6656
rect 5356 6604 5408 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 4610 6502 4662 6554
rect 4674 6502 4726 6554
rect 4738 6502 4790 6554
rect 4802 6502 4854 6554
rect 4866 6502 4918 6554
rect 6610 6502 6662 6554
rect 6674 6502 6726 6554
rect 6738 6502 6790 6554
rect 6802 6502 6854 6554
rect 6866 6502 6918 6554
rect 8610 6502 8662 6554
rect 8674 6502 8726 6554
rect 8738 6502 8790 6554
rect 8802 6502 8854 6554
rect 8866 6502 8918 6554
rect 2504 6400 2556 6452
rect 1584 6264 1636 6316
rect 1768 6264 1820 6316
rect 2228 6307 2280 6316
rect 2228 6273 2241 6307
rect 2241 6273 2275 6307
rect 2275 6273 2280 6307
rect 2228 6264 2280 6273
rect 2964 6264 3016 6316
rect 4160 6264 4212 6316
rect 1768 6128 1820 6180
rect 1860 6128 1912 6180
rect 3700 6239 3752 6248
rect 3700 6205 3709 6239
rect 3709 6205 3743 6239
rect 3743 6205 3752 6239
rect 3700 6196 3752 6205
rect 3884 6196 3936 6248
rect 4436 6264 4488 6316
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 5356 6400 5408 6452
rect 7104 6332 7156 6384
rect 7840 6332 7892 6384
rect 7472 6264 7524 6316
rect 8484 6264 8536 6316
rect 3424 6060 3476 6112
rect 4160 6060 4212 6112
rect 5448 6060 5500 6112
rect 6276 6060 6328 6112
rect 6736 6060 6788 6112
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 3950 5958 4002 6010
rect 4014 5958 4066 6010
rect 4078 5958 4130 6010
rect 4142 5958 4194 6010
rect 4206 5958 4258 6010
rect 5950 5958 6002 6010
rect 6014 5958 6066 6010
rect 6078 5958 6130 6010
rect 6142 5958 6194 6010
rect 6206 5958 6258 6010
rect 7950 5958 8002 6010
rect 8014 5958 8066 6010
rect 8078 5958 8130 6010
rect 8142 5958 8194 6010
rect 8206 5958 8258 6010
rect 1492 5856 1544 5908
rect 1860 5856 1912 5908
rect 7012 5856 7064 5908
rect 5172 5788 5224 5840
rect 5448 5720 5500 5772
rect 5816 5720 5868 5772
rect 1860 5584 1912 5636
rect 4436 5584 4488 5636
rect 6276 5695 6328 5704
rect 6276 5661 6283 5695
rect 6283 5661 6328 5695
rect 1768 5516 1820 5568
rect 5448 5516 5500 5568
rect 6276 5652 6328 5661
rect 7472 5788 7524 5840
rect 6368 5627 6420 5636
rect 6368 5593 6377 5627
rect 6377 5593 6411 5627
rect 6411 5593 6420 5627
rect 6368 5584 6420 5593
rect 6736 5652 6788 5704
rect 7840 5652 7892 5704
rect 8484 5652 8536 5704
rect 7380 5559 7432 5568
rect 7380 5525 7389 5559
rect 7389 5525 7423 5559
rect 7423 5525 7432 5559
rect 7380 5516 7432 5525
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 4610 5414 4662 5466
rect 4674 5414 4726 5466
rect 4738 5414 4790 5466
rect 4802 5414 4854 5466
rect 4866 5414 4918 5466
rect 6610 5414 6662 5466
rect 6674 5414 6726 5466
rect 6738 5414 6790 5466
rect 6802 5414 6854 5466
rect 6866 5414 6918 5466
rect 8610 5414 8662 5466
rect 8674 5414 8726 5466
rect 8738 5414 8790 5466
rect 8802 5414 8854 5466
rect 8866 5414 8918 5466
rect 2780 5312 2832 5364
rect 3332 5312 3384 5364
rect 3792 5312 3844 5364
rect 6368 5312 6420 5364
rect 940 5244 992 5296
rect 3424 5244 3476 5296
rect 3608 5176 3660 5228
rect 5080 5219 5132 5228
rect 5080 5185 5089 5219
rect 5089 5185 5123 5219
rect 5123 5185 5132 5219
rect 5080 5176 5132 5185
rect 5816 5176 5868 5228
rect 3240 5040 3292 5092
rect 4804 5015 4856 5024
rect 4804 4981 4813 5015
rect 4813 4981 4847 5015
rect 4847 4981 4856 5015
rect 4804 4972 4856 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 3950 4870 4002 4922
rect 4014 4870 4066 4922
rect 4078 4870 4130 4922
rect 4142 4870 4194 4922
rect 4206 4870 4258 4922
rect 5950 4870 6002 4922
rect 6014 4870 6066 4922
rect 6078 4870 6130 4922
rect 6142 4870 6194 4922
rect 6206 4870 6258 4922
rect 7950 4870 8002 4922
rect 8014 4870 8066 4922
rect 8078 4870 8130 4922
rect 8142 4870 8194 4922
rect 8206 4870 8258 4922
rect 1492 4768 1544 4820
rect 1676 4768 1728 4820
rect 2412 4768 2464 4820
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 5080 4768 5132 4820
rect 4528 4700 4580 4752
rect 4896 4700 4948 4752
rect 2412 4564 2464 4616
rect 2780 4539 2832 4548
rect 2780 4505 2789 4539
rect 2789 4505 2823 4539
rect 2823 4505 2832 4539
rect 3056 4564 3108 4616
rect 3332 4607 3384 4616
rect 3332 4573 3341 4607
rect 3341 4573 3375 4607
rect 3375 4573 3384 4607
rect 3332 4564 3384 4573
rect 4804 4564 4856 4616
rect 5632 4564 5684 4616
rect 5908 4564 5960 4616
rect 2780 4496 2832 4505
rect 3792 4539 3844 4548
rect 3792 4505 3801 4539
rect 3801 4505 3835 4539
rect 3835 4505 3844 4539
rect 3792 4496 3844 4505
rect 2136 4471 2188 4480
rect 2136 4437 2145 4471
rect 2145 4437 2179 4471
rect 2179 4437 2188 4471
rect 2136 4428 2188 4437
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 4896 4539 4948 4548
rect 4896 4505 4905 4539
rect 4905 4505 4939 4539
rect 4939 4505 4948 4539
rect 4896 4496 4948 4505
rect 6368 4428 6420 4480
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 4610 4326 4662 4378
rect 4674 4326 4726 4378
rect 4738 4326 4790 4378
rect 4802 4326 4854 4378
rect 4866 4326 4918 4378
rect 6610 4326 6662 4378
rect 6674 4326 6726 4378
rect 6738 4326 6790 4378
rect 6802 4326 6854 4378
rect 6866 4326 6918 4378
rect 8610 4326 8662 4378
rect 8674 4326 8726 4378
rect 8738 4326 8790 4378
rect 8802 4326 8854 4378
rect 8866 4326 8918 4378
rect 3792 4224 3844 4276
rect 4160 4224 4212 4276
rect 5448 4224 5500 4276
rect 2136 4156 2188 4208
rect 5172 4156 5224 4208
rect 5908 4199 5960 4208
rect 5908 4165 5917 4199
rect 5917 4165 5951 4199
rect 5951 4165 5960 4199
rect 5908 4156 5960 4165
rect 3056 4131 3108 4140
rect 3056 4097 3065 4131
rect 3065 4097 3099 4131
rect 3099 4097 3108 4131
rect 3056 4088 3108 4097
rect 3240 4020 3292 4072
rect 4896 4020 4948 4072
rect 5080 4020 5132 4072
rect 3424 3927 3476 3936
rect 3424 3893 3433 3927
rect 3433 3893 3467 3927
rect 3467 3893 3476 3927
rect 3424 3884 3476 3893
rect 5448 4131 5500 4140
rect 5448 4097 5457 4131
rect 5457 4097 5491 4131
rect 5491 4097 5500 4131
rect 5448 4088 5500 4097
rect 6460 4156 6512 4208
rect 5540 3952 5592 4004
rect 6276 4020 6328 4072
rect 7380 4131 7432 4140
rect 7380 4097 7389 4131
rect 7389 4097 7423 4131
rect 7423 4097 7432 4131
rect 7380 4088 7432 4097
rect 7564 4131 7616 4140
rect 7564 4097 7573 4131
rect 7573 4097 7607 4131
rect 7607 4097 7616 4131
rect 7564 4088 7616 4097
rect 5724 3884 5776 3936
rect 6000 3884 6052 3936
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 7012 3927 7064 3936
rect 7012 3893 7021 3927
rect 7021 3893 7055 3927
rect 7055 3893 7064 3927
rect 7012 3884 7064 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 3950 3782 4002 3834
rect 4014 3782 4066 3834
rect 4078 3782 4130 3834
rect 4142 3782 4194 3834
rect 4206 3782 4258 3834
rect 5950 3782 6002 3834
rect 6014 3782 6066 3834
rect 6078 3782 6130 3834
rect 6142 3782 6194 3834
rect 6206 3782 6258 3834
rect 7950 3782 8002 3834
rect 8014 3782 8066 3834
rect 8078 3782 8130 3834
rect 8142 3782 8194 3834
rect 8206 3782 8258 3834
rect 4528 3612 4580 3664
rect 6092 3680 6144 3732
rect 7564 3680 7616 3732
rect 4896 3544 4948 3596
rect 5540 3476 5592 3528
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 5816 3408 5868 3460
rect 6368 3544 6420 3596
rect 6736 3544 6788 3596
rect 9220 3476 9272 3528
rect 5724 3340 5776 3392
rect 6276 3383 6328 3392
rect 6276 3349 6285 3383
rect 6285 3349 6319 3383
rect 6319 3349 6328 3383
rect 6276 3340 6328 3349
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 4610 3238 4662 3290
rect 4674 3238 4726 3290
rect 4738 3238 4790 3290
rect 4802 3238 4854 3290
rect 4866 3238 4918 3290
rect 6610 3238 6662 3290
rect 6674 3238 6726 3290
rect 6738 3238 6790 3290
rect 6802 3238 6854 3290
rect 6866 3238 6918 3290
rect 8610 3238 8662 3290
rect 8674 3238 8726 3290
rect 8738 3238 8790 3290
rect 8802 3238 8854 3290
rect 8866 3238 8918 3290
rect 4528 3136 4580 3188
rect 5080 3136 5132 3188
rect 5172 3179 5224 3188
rect 5172 3145 5197 3179
rect 5197 3145 5224 3179
rect 5172 3136 5224 3145
rect 5632 3136 5684 3188
rect 5816 3179 5868 3188
rect 5816 3145 5825 3179
rect 5825 3145 5859 3179
rect 5859 3145 5868 3179
rect 5816 3136 5868 3145
rect 6092 3136 6144 3188
rect 6184 3179 6236 3188
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 7380 3136 7432 3188
rect 3148 3068 3200 3120
rect 2872 3000 2924 3052
rect 940 2796 992 2848
rect 6276 3000 6328 3052
rect 7012 3000 7064 3052
rect 7196 2864 7248 2916
rect 6460 2839 6512 2848
rect 6460 2805 6469 2839
rect 6469 2805 6503 2839
rect 6503 2805 6512 2839
rect 6460 2796 6512 2805
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 3950 2694 4002 2746
rect 4014 2694 4066 2746
rect 4078 2694 4130 2746
rect 4142 2694 4194 2746
rect 4206 2694 4258 2746
rect 5950 2694 6002 2746
rect 6014 2694 6066 2746
rect 6078 2694 6130 2746
rect 6142 2694 6194 2746
rect 6206 2694 6258 2746
rect 7950 2694 8002 2746
rect 8014 2694 8066 2746
rect 8078 2694 8130 2746
rect 8142 2694 8194 2746
rect 8206 2694 8258 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 2872 2635 2924 2644
rect 2872 2601 2881 2635
rect 2881 2601 2915 2635
rect 2915 2601 2924 2635
rect 2872 2592 2924 2601
rect 7196 2592 7248 2644
rect 8484 2592 8536 2644
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 6460 2388 6512 2440
rect 20 2320 72 2372
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 5172 2295 5224 2304
rect 5172 2261 5181 2295
rect 5181 2261 5215 2295
rect 5215 2261 5224 2295
rect 5172 2252 5224 2261
rect 9036 2252 9088 2304
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
rect 4610 2150 4662 2202
rect 4674 2150 4726 2202
rect 4738 2150 4790 2202
rect 4802 2150 4854 2202
rect 4866 2150 4918 2202
rect 6610 2150 6662 2202
rect 6674 2150 6726 2202
rect 6738 2150 6790 2202
rect 6802 2150 6854 2202
rect 6866 2150 6918 2202
rect 8610 2150 8662 2202
rect 8674 2150 8726 2202
rect 8738 2150 8790 2202
rect 8802 2150 8854 2202
rect 8866 2150 8918 2202
<< metal2 >>
rect 1306 11618 1362 12418
rect 4526 11618 4582 12418
rect 7102 11778 7158 12418
rect 7102 11750 7420 11778
rect 7102 11618 7158 11750
rect 1320 9654 1348 11618
rect 1858 11384 1914 11393
rect 1858 11319 1914 11328
rect 1872 9654 1900 11319
rect 2610 9820 2918 9829
rect 2610 9818 2616 9820
rect 2672 9818 2696 9820
rect 2752 9818 2776 9820
rect 2832 9818 2856 9820
rect 2912 9818 2918 9820
rect 2672 9766 2674 9818
rect 2854 9766 2856 9818
rect 2610 9764 2616 9766
rect 2672 9764 2696 9766
rect 2752 9764 2776 9766
rect 2832 9764 2856 9766
rect 2912 9764 2918 9766
rect 2610 9755 2918 9764
rect 4540 9654 4568 11618
rect 4610 9820 4918 9829
rect 4610 9818 4616 9820
rect 4672 9818 4696 9820
rect 4752 9818 4776 9820
rect 4832 9818 4856 9820
rect 4912 9818 4918 9820
rect 4672 9766 4674 9818
rect 4854 9766 4856 9818
rect 4610 9764 4616 9766
rect 4672 9764 4696 9766
rect 4752 9764 4776 9766
rect 4832 9764 4856 9766
rect 4912 9764 4918 9766
rect 4610 9755 4918 9764
rect 6610 9820 6918 9829
rect 6610 9818 6616 9820
rect 6672 9818 6696 9820
rect 6752 9818 6776 9820
rect 6832 9818 6856 9820
rect 6912 9818 6918 9820
rect 6672 9766 6674 9818
rect 6854 9766 6856 9818
rect 6610 9764 6616 9766
rect 6672 9764 6696 9766
rect 6752 9764 6776 9766
rect 6832 9764 6856 9766
rect 6912 9764 6918 9766
rect 6610 9755 6918 9764
rect 7392 9654 7420 11750
rect 9678 11618 9734 12418
rect 8610 9820 8918 9829
rect 8610 9818 8616 9820
rect 8672 9818 8696 9820
rect 8752 9818 8776 9820
rect 8832 9818 8856 9820
rect 8912 9818 8918 9820
rect 8672 9766 8674 9818
rect 8854 9766 8856 9818
rect 8610 9764 8616 9766
rect 8672 9764 8696 9766
rect 8752 9764 8776 9766
rect 8832 9764 8856 9766
rect 8912 9764 8918 9766
rect 8610 9755 8918 9764
rect 9692 9654 9720 11618
rect 1308 9648 1360 9654
rect 1308 9590 1360 9596
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7748 9648 7800 9654
rect 9680 9648 9732 9654
rect 7748 9590 7800 9596
rect 8942 9616 8998 9625
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 1504 8906 1532 9318
rect 938 8871 994 8880
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1504 5914 1532 8842
rect 1688 7954 1716 9318
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 3950 9276 4258 9285
rect 3950 9274 3956 9276
rect 4012 9274 4036 9276
rect 4092 9274 4116 9276
rect 4172 9274 4196 9276
rect 4252 9274 4258 9276
rect 4012 9222 4014 9274
rect 4194 9222 4196 9274
rect 3950 9220 3956 9222
rect 4012 9220 4036 9222
rect 4092 9220 4116 9222
rect 4172 9220 4196 9222
rect 4252 9220 4258 9222
rect 3950 9211 4258 9220
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1676 7948 1728 7954
rect 1676 7890 1728 7896
rect 1688 7274 1716 7890
rect 1676 7268 1728 7274
rect 1676 7210 1728 7216
rect 1780 6322 1808 8910
rect 3252 8894 3464 8922
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 3252 8634 3280 8894
rect 3436 8838 3464 8894
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 3344 8498 3372 8774
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1860 7880 1912 7886
rect 1860 7822 1912 7828
rect 1872 7478 1900 7822
rect 2516 7698 2544 8434
rect 2976 8294 3004 8434
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2424 7670 2544 7698
rect 1860 7472 1912 7478
rect 1860 7414 1912 7420
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 1584 6316 1636 6322
rect 1768 6316 1820 6322
rect 1584 6258 1636 6264
rect 1688 6276 1768 6304
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 938 5536 994 5545
rect 938 5471 994 5480
rect 952 5302 980 5471
rect 940 5296 992 5302
rect 940 5238 992 5244
rect 1504 4826 1532 5850
rect 1492 4820 1544 4826
rect 1492 4762 1544 4768
rect 940 2848 992 2854
rect 938 2816 940 2825
rect 992 2816 994 2825
rect 938 2751 994 2760
rect 1596 2650 1624 6258
rect 1688 4826 1716 6276
rect 1768 6258 1820 6264
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2240 6202 2268 6258
rect 2424 6202 2452 7670
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2504 7472 2556 7478
rect 2504 7414 2556 7420
rect 2516 6458 2544 7414
rect 2964 7268 3016 7274
rect 2964 7210 3016 7216
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2976 6322 3004 7210
rect 2964 6316 3016 6322
rect 2964 6258 3016 6264
rect 1768 6180 1820 6186
rect 1768 6122 1820 6128
rect 1860 6180 1912 6186
rect 2240 6174 2452 6202
rect 1860 6122 1912 6128
rect 1780 5574 1808 6122
rect 1872 5914 1900 6122
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 1676 4820 1728 4826
rect 1676 4762 1728 4768
rect 1872 4622 1900 5578
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2332 4706 2360 6174
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 2412 4820 2464 4826
rect 2412 4762 2464 4768
rect 2148 4678 2360 4706
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 2148 4486 2176 4678
rect 2424 4622 2452 4762
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2792 4554 2820 5306
rect 3056 4616 3108 4622
rect 3056 4558 3108 4564
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2148 4214 2176 4422
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 2136 4208 2188 4214
rect 2136 4150 2188 4156
rect 3068 4146 3096 4558
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 1950 3771 2258 3780
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 3160 3126 3188 8298
rect 3528 8294 3556 8978
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3620 8634 3648 8774
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3712 8514 3740 8774
rect 3620 8486 3740 8514
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3240 5092 3292 5098
rect 3240 5034 3292 5040
rect 3252 4078 3280 5034
rect 3344 4622 3372 5306
rect 3436 5302 3464 6054
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 3620 5234 3648 8486
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3712 6254 3740 8298
rect 3700 6248 3752 6254
rect 3700 6190 3752 6196
rect 3804 5370 3832 8502
rect 4172 8498 4200 8910
rect 4610 8732 4918 8741
rect 4610 8730 4616 8732
rect 4672 8730 4696 8732
rect 4752 8730 4776 8732
rect 4832 8730 4856 8732
rect 4912 8730 4918 8732
rect 4672 8678 4674 8730
rect 4854 8678 4856 8730
rect 4610 8676 4616 8678
rect 4672 8676 4696 8678
rect 4752 8676 4776 8678
rect 4832 8676 4856 8678
rect 4912 8676 4918 8678
rect 4610 8667 4918 8676
rect 5000 8634 5028 9318
rect 5950 9276 6258 9285
rect 5950 9274 5956 9276
rect 6012 9274 6036 9276
rect 6092 9274 6116 9276
rect 6172 9274 6196 9276
rect 6252 9274 6258 9276
rect 6012 9222 6014 9274
rect 6194 9222 6196 9274
rect 5950 9220 5956 9222
rect 6012 9220 6036 9222
rect 6092 9220 6116 9222
rect 6172 9220 6196 9222
rect 6252 9220 6258 9222
rect 5950 9211 6258 9220
rect 7300 9178 7328 9522
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 3950 8188 4258 8197
rect 3950 8186 3956 8188
rect 4012 8186 4036 8188
rect 4092 8186 4116 8188
rect 4172 8186 4196 8188
rect 4252 8186 4258 8188
rect 4012 8134 4014 8186
rect 4194 8134 4196 8186
rect 3950 8132 3956 8134
rect 4012 8132 4036 8134
rect 4092 8132 4116 8134
rect 4172 8132 4196 8134
rect 4252 8132 4258 8134
rect 3950 8123 4258 8132
rect 4610 7644 4918 7653
rect 4610 7642 4616 7644
rect 4672 7642 4696 7644
rect 4752 7642 4776 7644
rect 4832 7642 4856 7644
rect 4912 7642 4918 7644
rect 4672 7590 4674 7642
rect 4854 7590 4856 7642
rect 4610 7588 4616 7590
rect 4672 7588 4696 7590
rect 4752 7588 4776 7590
rect 4832 7588 4856 7590
rect 4912 7588 4918 7590
rect 4610 7579 4918 7588
rect 5000 7274 5028 8230
rect 5184 7954 5212 8230
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5080 7880 5132 7886
rect 5080 7822 5132 7828
rect 5092 7546 5120 7822
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7410 5212 7890
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 7410 5396 7686
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 3950 7100 4258 7109
rect 3950 7098 3956 7100
rect 4012 7098 4036 7100
rect 4092 7098 4116 7100
rect 4172 7098 4196 7100
rect 4252 7098 4258 7100
rect 4012 7046 4014 7098
rect 4194 7046 4196 7098
rect 3950 7044 3956 7046
rect 4012 7044 4036 7046
rect 4092 7044 4116 7046
rect 4172 7044 4196 7046
rect 4252 7044 4258 7046
rect 3950 7035 4258 7044
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4172 6322 4200 6598
rect 4540 6322 4568 7142
rect 5368 6662 5396 7346
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 4610 6556 4918 6565
rect 4610 6554 4616 6556
rect 4672 6554 4696 6556
rect 4752 6554 4776 6556
rect 4832 6554 4856 6556
rect 4912 6554 4918 6556
rect 4672 6502 4674 6554
rect 4854 6502 4856 6554
rect 4610 6500 4616 6502
rect 4672 6500 4696 6502
rect 4752 6500 4776 6502
rect 4832 6500 4856 6502
rect 4912 6500 4918 6502
rect 4610 6491 4918 6500
rect 5368 6458 5396 6598
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4436 6316 4488 6322
rect 4436 6258 4488 6264
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 3884 6248 3936 6254
rect 3936 6196 4200 6202
rect 3884 6190 4200 6196
rect 3896 6174 4200 6190
rect 4172 6118 4200 6174
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 3950 6012 4258 6021
rect 3950 6010 3956 6012
rect 4012 6010 4036 6012
rect 4092 6010 4116 6012
rect 4172 6010 4196 6012
rect 4252 6010 4258 6012
rect 4012 5958 4014 6010
rect 4194 5958 4196 6010
rect 3950 5956 3956 5958
rect 4012 5956 4036 5958
rect 4092 5956 4116 5958
rect 4172 5956 4196 5958
rect 4252 5956 4258 5958
rect 3950 5947 4258 5956
rect 4448 5642 4476 6258
rect 5448 6112 5500 6118
rect 5448 6054 5500 6060
rect 5172 5840 5224 5846
rect 5172 5782 5224 5788
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4610 5468 4918 5477
rect 4610 5466 4616 5468
rect 4672 5466 4696 5468
rect 4752 5466 4776 5468
rect 4832 5466 4856 5468
rect 4912 5466 4918 5468
rect 4672 5414 4674 5466
rect 4854 5414 4856 5466
rect 4610 5412 4616 5414
rect 4672 5412 4696 5414
rect 4752 5412 4776 5414
rect 4832 5412 4856 5414
rect 4912 5412 4918 5414
rect 4610 5403 4918 5412
rect 3792 5364 3844 5370
rect 3792 5306 3844 5312
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 3950 4924 4258 4933
rect 3950 4922 3956 4924
rect 4012 4922 4036 4924
rect 4092 4922 4116 4924
rect 4172 4922 4196 4924
rect 4252 4922 4258 4924
rect 4012 4870 4014 4922
rect 4194 4870 4196 4922
rect 3950 4868 3956 4870
rect 4012 4868 4036 4870
rect 4092 4868 4116 4870
rect 4172 4868 4196 4870
rect 4252 4868 4258 4870
rect 3950 4859 4258 4868
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3436 3942 3464 4762
rect 4528 4752 4580 4758
rect 4528 4694 4580 4700
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3804 4282 3832 4490
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 4172 4282 4200 4422
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3950 3836 4258 3845
rect 3950 3834 3956 3836
rect 4012 3834 4036 3836
rect 4092 3834 4116 3836
rect 4172 3834 4196 3836
rect 4252 3834 4258 3836
rect 4012 3782 4014 3834
rect 4194 3782 4196 3834
rect 3950 3780 3956 3782
rect 4012 3780 4036 3782
rect 4092 3780 4116 3782
rect 4172 3780 4196 3782
rect 4252 3780 4258 3782
rect 3950 3771 4258 3780
rect 4540 3670 4568 4694
rect 4816 4622 4844 4966
rect 5092 4826 5120 5170
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 4896 4752 4948 4758
rect 4896 4694 4948 4700
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4908 4554 4936 4694
rect 4896 4548 4948 4554
rect 4896 4490 4948 4496
rect 4610 4380 4918 4389
rect 4610 4378 4616 4380
rect 4672 4378 4696 4380
rect 4752 4378 4776 4380
rect 4832 4378 4856 4380
rect 4912 4378 4918 4380
rect 4672 4326 4674 4378
rect 4854 4326 4856 4378
rect 4610 4324 4616 4326
rect 4672 4324 4696 4326
rect 4752 4324 4776 4326
rect 4832 4324 4856 4326
rect 4912 4324 4918 4326
rect 4610 4315 4918 4324
rect 5184 4214 5212 5782
rect 5460 5778 5488 6054
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5460 4282 5488 5510
rect 5644 4622 5672 7822
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5448 4276 5500 4282
rect 5448 4218 5500 4224
rect 5172 4208 5224 4214
rect 5644 4162 5672 4558
rect 5172 4150 5224 4156
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 5080 4072 5132 4078
rect 5080 4014 5132 4020
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4540 3194 4568 3606
rect 4908 3602 4936 4014
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 4610 3292 4918 3301
rect 4610 3290 4616 3292
rect 4672 3290 4696 3292
rect 4752 3290 4776 3292
rect 4832 3290 4856 3292
rect 4912 3290 4918 3292
rect 4672 3238 4674 3290
rect 4854 3238 4856 3290
rect 4610 3236 4616 3238
rect 4672 3236 4696 3238
rect 4752 3236 4776 3238
rect 4832 3236 4856 3238
rect 4912 3236 4918 3238
rect 4610 3227 4918 3236
rect 5092 3194 5120 4014
rect 5184 3194 5212 4150
rect 5460 4146 5672 4162
rect 5448 4140 5672 4146
rect 5500 4134 5672 4140
rect 5736 4162 5764 8910
rect 6610 8732 6918 8741
rect 6610 8730 6616 8732
rect 6672 8730 6696 8732
rect 6752 8730 6776 8732
rect 6832 8730 6856 8732
rect 6912 8730 6918 8732
rect 6672 8678 6674 8730
rect 6854 8678 6856 8730
rect 6610 8676 6616 8678
rect 6672 8676 6696 8678
rect 6752 8676 6776 8678
rect 6832 8676 6856 8678
rect 6912 8676 6918 8678
rect 6610 8667 6918 8676
rect 5950 8188 6258 8197
rect 5950 8186 5956 8188
rect 6012 8186 6036 8188
rect 6092 8186 6116 8188
rect 6172 8186 6196 8188
rect 6252 8186 6258 8188
rect 6012 8134 6014 8186
rect 6194 8134 6196 8186
rect 5950 8132 5956 8134
rect 6012 8132 6036 8134
rect 6092 8132 6116 8134
rect 6172 8132 6196 8134
rect 6252 8132 6258 8134
rect 5950 8123 6258 8132
rect 7760 8090 7788 9590
rect 9680 9590 9732 9596
rect 8942 9551 8944 9560
rect 8996 9551 8998 9560
rect 8944 9522 8996 9528
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 5920 7750 5948 7822
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5828 7546 5856 7686
rect 6472 7546 6500 7822
rect 6610 7644 6918 7653
rect 6610 7642 6616 7644
rect 6672 7642 6696 7644
rect 6752 7642 6776 7644
rect 6832 7642 6856 7644
rect 6912 7642 6918 7644
rect 6672 7590 6674 7642
rect 6854 7590 6856 7642
rect 6610 7588 6616 7590
rect 6672 7588 6696 7590
rect 6752 7588 6776 7590
rect 6832 7588 6856 7590
rect 6912 7588 6918 7590
rect 6610 7579 6918 7588
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 5950 7100 6258 7109
rect 5950 7098 5956 7100
rect 6012 7098 6036 7100
rect 6092 7098 6116 7100
rect 6172 7098 6196 7100
rect 6252 7098 6258 7100
rect 6012 7046 6014 7098
rect 6194 7046 6196 7098
rect 5950 7044 5956 7046
rect 6012 7044 6036 7046
rect 6092 7044 6116 7046
rect 6172 7044 6196 7046
rect 6252 7044 6258 7046
rect 5950 7035 6258 7044
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 5950 6012 6258 6021
rect 5950 6010 5956 6012
rect 6012 6010 6036 6012
rect 6092 6010 6116 6012
rect 6172 6010 6196 6012
rect 6252 6010 6258 6012
rect 6012 5958 6014 6010
rect 6194 5958 6196 6010
rect 5950 5956 5956 5958
rect 6012 5956 6036 5958
rect 6092 5956 6116 5958
rect 6172 5956 6196 5958
rect 6252 5956 6258 5958
rect 5950 5947 6258 5956
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5828 5234 5856 5714
rect 6288 5710 6316 6054
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6380 5370 6408 5578
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5950 4924 6258 4933
rect 5950 4922 5956 4924
rect 6012 4922 6036 4924
rect 6092 4922 6116 4924
rect 6172 4922 6196 4924
rect 6252 4922 6258 4924
rect 6012 4870 6014 4922
rect 6194 4870 6196 4922
rect 5950 4868 5956 4870
rect 6012 4868 6036 4870
rect 6092 4868 6116 4870
rect 6172 4868 6196 4870
rect 6252 4868 6258 4870
rect 5950 4859 6258 4868
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5920 4214 5948 4558
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 5908 4208 5960 4214
rect 5736 4134 5856 4162
rect 5908 4150 5960 4156
rect 5448 4082 5500 4088
rect 5828 4026 5856 4134
rect 6276 4072 6328 4078
rect 5540 4004 5592 4010
rect 5828 3998 6040 4026
rect 6276 4014 6328 4020
rect 5540 3946 5592 3952
rect 5552 3534 5580 3946
rect 6012 3942 6040 3998
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 5644 3194 5672 3470
rect 5736 3398 5764 3878
rect 5950 3836 6258 3845
rect 5950 3834 5956 3836
rect 6012 3834 6036 3836
rect 6092 3834 6116 3836
rect 6172 3834 6196 3836
rect 6252 3834 6258 3836
rect 6012 3782 6014 3834
rect 6194 3782 6196 3834
rect 5950 3780 5956 3782
rect 6012 3780 6036 3782
rect 6092 3780 6116 3782
rect 6172 3780 6196 3782
rect 6252 3780 6258 3782
rect 5950 3771 6258 3780
rect 6092 3732 6144 3738
rect 6092 3674 6144 3680
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5828 3194 5856 3402
rect 6104 3194 6132 3674
rect 6288 3618 6316 4014
rect 6196 3590 6316 3618
rect 6380 3602 6408 4422
rect 6472 4214 6500 7142
rect 6610 6556 6918 6565
rect 6610 6554 6616 6556
rect 6672 6554 6696 6556
rect 6752 6554 6776 6556
rect 6832 6554 6856 6556
rect 6912 6554 6918 6556
rect 6672 6502 6674 6554
rect 6854 6502 6856 6554
rect 6610 6500 6616 6502
rect 6672 6500 6696 6502
rect 6752 6500 6776 6502
rect 6832 6500 6856 6502
rect 6912 6500 6918 6502
rect 6610 6491 6918 6500
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6748 5710 6776 6054
rect 7024 5914 7052 7822
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7410 7144 7686
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 7116 6390 7144 7346
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7300 7002 7328 7278
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7852 6866 7880 9318
rect 7950 9276 8258 9285
rect 7950 9274 7956 9276
rect 8012 9274 8036 9276
rect 8092 9274 8116 9276
rect 8172 9274 8196 9276
rect 8252 9274 8258 9276
rect 8012 9222 8014 9274
rect 8194 9222 8196 9274
rect 7950 9220 7956 9222
rect 8012 9220 8036 9222
rect 8092 9220 8116 9222
rect 8172 9220 8196 9222
rect 8252 9220 8258 9222
rect 7950 9211 8258 9220
rect 8610 8732 8918 8741
rect 8610 8730 8616 8732
rect 8672 8730 8696 8732
rect 8752 8730 8776 8732
rect 8832 8730 8856 8732
rect 8912 8730 8918 8732
rect 8672 8678 8674 8730
rect 8854 8678 8856 8730
rect 8610 8676 8616 8678
rect 8672 8676 8696 8678
rect 8752 8676 8776 8678
rect 8832 8676 8856 8678
rect 8912 8676 8918 8678
rect 8610 8667 8918 8676
rect 7950 8188 8258 8197
rect 7950 8186 7956 8188
rect 8012 8186 8036 8188
rect 8092 8186 8116 8188
rect 8172 8186 8196 8188
rect 8252 8186 8258 8188
rect 8012 8134 8014 8186
rect 8194 8134 8196 8186
rect 7950 8132 7956 8134
rect 8012 8132 8036 8134
rect 8092 8132 8116 8134
rect 8172 8132 8196 8134
rect 8252 8132 8258 8134
rect 7950 8123 8258 8132
rect 8610 7644 8918 7653
rect 8610 7642 8616 7644
rect 8672 7642 8696 7644
rect 8752 7642 8776 7644
rect 8832 7642 8856 7644
rect 8912 7642 8918 7644
rect 8672 7590 8674 7642
rect 8854 7590 8856 7642
rect 8610 7588 8616 7590
rect 8672 7588 8696 7590
rect 8752 7588 8776 7590
rect 8832 7588 8856 7590
rect 8912 7588 8918 7590
rect 8610 7579 8918 7588
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 7950 7100 8258 7109
rect 7950 7098 7956 7100
rect 8012 7098 8036 7100
rect 8092 7098 8116 7100
rect 8172 7098 8196 7100
rect 8252 7098 8258 7100
rect 8012 7046 8014 7098
rect 8194 7046 8196 7098
rect 7950 7044 7956 7046
rect 8012 7044 8036 7046
rect 8092 7044 8116 7046
rect 8172 7044 8196 7046
rect 8252 7044 8258 7046
rect 7950 7035 8258 7044
rect 9232 6905 9260 7278
rect 9218 6896 9274 6905
rect 7840 6860 7892 6866
rect 9218 6831 9274 6840
rect 7840 6802 7892 6808
rect 7852 6390 7880 6802
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 7484 5846 7512 6258
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7852 5710 7880 6326
rect 8496 6322 8524 6666
rect 8610 6556 8918 6565
rect 8610 6554 8616 6556
rect 8672 6554 8696 6556
rect 8752 6554 8776 6556
rect 8832 6554 8856 6556
rect 8912 6554 8918 6556
rect 8672 6502 8674 6554
rect 8854 6502 8856 6554
rect 8610 6500 8616 6502
rect 8672 6500 8696 6502
rect 8752 6500 8776 6502
rect 8832 6500 8856 6502
rect 8912 6500 8918 6502
rect 8610 6491 8918 6500
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 7950 6012 8258 6021
rect 7950 6010 7956 6012
rect 8012 6010 8036 6012
rect 8092 6010 8116 6012
rect 8172 6010 8196 6012
rect 8252 6010 8258 6012
rect 8012 5958 8014 6010
rect 8194 5958 8196 6010
rect 7950 5956 7956 5958
rect 8012 5956 8036 5958
rect 8092 5956 8116 5958
rect 8172 5956 8196 5958
rect 8252 5956 8258 5958
rect 7950 5947 8258 5956
rect 8496 5710 8524 6258
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 8484 5704 8536 5710
rect 8484 5646 8536 5652
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 6610 5468 6918 5477
rect 6610 5466 6616 5468
rect 6672 5466 6696 5468
rect 6752 5466 6776 5468
rect 6832 5466 6856 5468
rect 6912 5466 6918 5468
rect 6672 5414 6674 5466
rect 6854 5414 6856 5466
rect 6610 5412 6616 5414
rect 6672 5412 6696 5414
rect 6752 5412 6776 5414
rect 6832 5412 6856 5414
rect 6912 5412 6918 5414
rect 6610 5403 6918 5412
rect 6610 4380 6918 4389
rect 6610 4378 6616 4380
rect 6672 4378 6696 4380
rect 6752 4378 6776 4380
rect 6832 4378 6856 4380
rect 6912 4378 6918 4380
rect 6672 4326 6674 4378
rect 6854 4326 6856 4378
rect 6610 4324 6616 4326
rect 6672 4324 6696 4326
rect 6752 4324 6776 4326
rect 6832 4324 6856 4326
rect 6912 4324 6918 4326
rect 6610 4315 6918 4324
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 7392 4146 7420 5510
rect 7950 4924 8258 4933
rect 7950 4922 7956 4924
rect 8012 4922 8036 4924
rect 8092 4922 8116 4924
rect 8172 4922 8196 4924
rect 8252 4922 8258 4924
rect 8012 4870 8014 4922
rect 8194 4870 8196 4922
rect 7950 4868 7956 4870
rect 8012 4868 8036 4870
rect 8092 4868 8116 4870
rect 8172 4868 8196 4870
rect 8252 4868 8258 4870
rect 7950 4859 8258 4868
rect 7380 4140 7432 4146
rect 7380 4082 7432 4088
rect 7564 4140 7616 4146
rect 7564 4082 7616 4088
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6748 3602 6776 3878
rect 6368 3596 6420 3602
rect 6196 3194 6224 3590
rect 6368 3538 6420 3544
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5816 3188 5868 3194
rect 5816 3130 5868 3136
rect 6092 3188 6144 3194
rect 6092 3130 6144 3136
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 6288 3058 6316 3334
rect 6610 3292 6918 3301
rect 6610 3290 6616 3292
rect 6672 3290 6696 3292
rect 6752 3290 6776 3292
rect 6832 3290 6856 3292
rect 6912 3290 6918 3292
rect 6672 3238 6674 3290
rect 6854 3238 6856 3290
rect 6610 3236 6616 3238
rect 6672 3236 6696 3238
rect 6752 3236 6776 3238
rect 6832 3236 6856 3238
rect 6912 3236 6918 3238
rect 6610 3227 6918 3236
rect 7024 3058 7052 3878
rect 7392 3194 7420 4082
rect 7576 3738 7604 4082
rect 7950 3836 8258 3845
rect 7950 3834 7956 3836
rect 8012 3834 8036 3836
rect 8092 3834 8116 3836
rect 8172 3834 8196 3836
rect 8252 3834 8258 3836
rect 8012 3782 8014 3834
rect 8194 3782 8196 3834
rect 7950 3780 7956 3782
rect 8012 3780 8036 3782
rect 8092 3780 8116 3782
rect 8172 3780 8196 3782
rect 8252 3780 8258 3782
rect 7950 3771 8258 3780
rect 7564 3732 7616 3738
rect 7564 3674 7616 3680
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2884 2650 2912 2994
rect 7196 2916 7248 2922
rect 7196 2858 7248 2864
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 3950 2748 4258 2757
rect 3950 2746 3956 2748
rect 4012 2746 4036 2748
rect 4092 2746 4116 2748
rect 4172 2746 4196 2748
rect 4252 2746 4258 2748
rect 4012 2694 4014 2746
rect 4194 2694 4196 2746
rect 3950 2692 3956 2694
rect 4012 2692 4036 2694
rect 4092 2692 4116 2694
rect 4172 2692 4196 2694
rect 4252 2692 4258 2694
rect 3950 2683 4258 2692
rect 5950 2748 6258 2757
rect 5950 2746 5956 2748
rect 6012 2746 6036 2748
rect 6092 2746 6116 2748
rect 6172 2746 6196 2748
rect 6252 2746 6258 2748
rect 6012 2694 6014 2746
rect 6194 2694 6196 2746
rect 5950 2692 5956 2694
rect 6012 2692 6036 2694
rect 6092 2692 6116 2694
rect 6172 2692 6196 2694
rect 6252 2692 6258 2694
rect 5950 2683 6258 2692
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 2872 2644 2924 2650
rect 2872 2586 2924 2592
rect 6472 2446 6500 2790
rect 7208 2650 7236 2858
rect 7950 2748 8258 2757
rect 7950 2746 7956 2748
rect 8012 2746 8036 2748
rect 8092 2746 8116 2748
rect 8172 2746 8196 2748
rect 8252 2746 8258 2748
rect 8012 2694 8014 2746
rect 8194 2694 8196 2746
rect 7950 2692 7956 2694
rect 8012 2692 8036 2694
rect 8092 2692 8116 2694
rect 8172 2692 8196 2694
rect 8252 2692 8258 2694
rect 7950 2683 8258 2692
rect 8496 2650 8524 5646
rect 8610 5468 8918 5477
rect 8610 5466 8616 5468
rect 8672 5466 8696 5468
rect 8752 5466 8776 5468
rect 8832 5466 8856 5468
rect 8912 5466 8918 5468
rect 8672 5414 8674 5466
rect 8854 5414 8856 5466
rect 8610 5412 8616 5414
rect 8672 5412 8696 5414
rect 8752 5412 8776 5414
rect 8832 5412 8856 5414
rect 8912 5412 8918 5414
rect 8610 5403 8918 5412
rect 8610 4380 8918 4389
rect 8610 4378 8616 4380
rect 8672 4378 8696 4380
rect 8752 4378 8776 4380
rect 8832 4378 8856 4380
rect 8912 4378 8918 4380
rect 8672 4326 8674 4378
rect 8854 4326 8856 4378
rect 8610 4324 8616 4326
rect 8672 4324 8696 4326
rect 8752 4324 8776 4326
rect 8832 4324 8856 4326
rect 8912 4324 8918 4326
rect 8610 4315 8918 4324
rect 9220 3528 9272 3534
rect 9218 3496 9220 3505
rect 9272 3496 9274 3505
rect 9218 3431 9274 3440
rect 8610 3292 8918 3301
rect 8610 3290 8616 3292
rect 8672 3290 8696 3292
rect 8752 3290 8776 3292
rect 8832 3290 8856 3292
rect 8912 3290 8918 3292
rect 8672 3238 8674 3290
rect 8854 3238 8856 3290
rect 8610 3236 8616 3238
rect 8672 3236 8696 3238
rect 8752 3236 8776 3238
rect 8832 3236 8856 3238
rect 8912 3236 8918 3238
rect 8610 3227 8918 3236
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 8484 2644 8536 2650
rect 8484 2586 8536 2592
rect 2688 2440 2740 2446
rect 2516 2388 2688 2394
rect 2516 2382 2740 2388
rect 6460 2440 6512 2446
rect 8484 2440 8536 2446
rect 6460 2382 6512 2388
rect 8404 2400 8484 2428
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 2516 2366 2728 2382
rect 32 800 60 2314
rect 2516 1306 2544 2366
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 2610 2204 2918 2213
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 4610 2204 4918 2213
rect 4610 2202 4616 2204
rect 4672 2202 4696 2204
rect 4752 2202 4776 2204
rect 4832 2202 4856 2204
rect 4912 2202 4918 2204
rect 4672 2150 4674 2202
rect 4854 2150 4856 2202
rect 4610 2148 4616 2150
rect 4672 2148 4696 2150
rect 4752 2148 4776 2150
rect 4832 2148 4856 2150
rect 4912 2148 4918 2150
rect 4610 2139 4918 2148
rect 2516 1278 2636 1306
rect 2608 800 2636 1278
rect 5184 800 5212 2246
rect 6610 2204 6918 2213
rect 6610 2202 6616 2204
rect 6672 2202 6696 2204
rect 6752 2202 6776 2204
rect 6832 2202 6856 2204
rect 6912 2202 6918 2204
rect 6672 2150 6674 2202
rect 6854 2150 6856 2202
rect 6610 2148 6616 2150
rect 6672 2148 6696 2150
rect 6752 2148 6776 2150
rect 6832 2148 6856 2150
rect 6912 2148 6918 2150
rect 6610 2139 6918 2148
rect 8404 800 8432 2400
rect 8484 2382 8536 2388
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 8610 2204 8918 2213
rect 8610 2202 8616 2204
rect 8672 2202 8696 2204
rect 8752 2202 8776 2204
rect 8832 2202 8856 2204
rect 8912 2202 8918 2204
rect 8672 2150 8674 2202
rect 8854 2150 8856 2202
rect 8610 2148 8616 2150
rect 8672 2148 8696 2150
rect 8752 2148 8776 2150
rect 8832 2148 8856 2150
rect 8912 2148 8918 2150
rect 8610 2139 8918 2148
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 8390 0 8446 800
rect 9048 785 9076 2246
rect 9034 776 9090 785
rect 9034 711 9090 720
<< via2 >>
rect 1858 11328 1914 11384
rect 2616 9818 2672 9820
rect 2696 9818 2752 9820
rect 2776 9818 2832 9820
rect 2856 9818 2912 9820
rect 2616 9766 2662 9818
rect 2662 9766 2672 9818
rect 2696 9766 2726 9818
rect 2726 9766 2738 9818
rect 2738 9766 2752 9818
rect 2776 9766 2790 9818
rect 2790 9766 2802 9818
rect 2802 9766 2832 9818
rect 2856 9766 2866 9818
rect 2866 9766 2912 9818
rect 2616 9764 2672 9766
rect 2696 9764 2752 9766
rect 2776 9764 2832 9766
rect 2856 9764 2912 9766
rect 4616 9818 4672 9820
rect 4696 9818 4752 9820
rect 4776 9818 4832 9820
rect 4856 9818 4912 9820
rect 4616 9766 4662 9818
rect 4662 9766 4672 9818
rect 4696 9766 4726 9818
rect 4726 9766 4738 9818
rect 4738 9766 4752 9818
rect 4776 9766 4790 9818
rect 4790 9766 4802 9818
rect 4802 9766 4832 9818
rect 4856 9766 4866 9818
rect 4866 9766 4912 9818
rect 4616 9764 4672 9766
rect 4696 9764 4752 9766
rect 4776 9764 4832 9766
rect 4856 9764 4912 9766
rect 6616 9818 6672 9820
rect 6696 9818 6752 9820
rect 6776 9818 6832 9820
rect 6856 9818 6912 9820
rect 6616 9766 6662 9818
rect 6662 9766 6672 9818
rect 6696 9766 6726 9818
rect 6726 9766 6738 9818
rect 6738 9766 6752 9818
rect 6776 9766 6790 9818
rect 6790 9766 6802 9818
rect 6802 9766 6832 9818
rect 6856 9766 6866 9818
rect 6866 9766 6912 9818
rect 6616 9764 6672 9766
rect 6696 9764 6752 9766
rect 6776 9764 6832 9766
rect 6856 9764 6912 9766
rect 8616 9818 8672 9820
rect 8696 9818 8752 9820
rect 8776 9818 8832 9820
rect 8856 9818 8912 9820
rect 8616 9766 8662 9818
rect 8662 9766 8672 9818
rect 8696 9766 8726 9818
rect 8726 9766 8738 9818
rect 8738 9766 8752 9818
rect 8776 9766 8790 9818
rect 8790 9766 8802 9818
rect 8802 9766 8832 9818
rect 8856 9766 8866 9818
rect 8866 9766 8912 9818
rect 8616 9764 8672 9766
rect 8696 9764 8752 9766
rect 8776 9764 8832 9766
rect 8856 9764 8912 9766
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 3956 9274 4012 9276
rect 4036 9274 4092 9276
rect 4116 9274 4172 9276
rect 4196 9274 4252 9276
rect 3956 9222 4002 9274
rect 4002 9222 4012 9274
rect 4036 9222 4066 9274
rect 4066 9222 4078 9274
rect 4078 9222 4092 9274
rect 4116 9222 4130 9274
rect 4130 9222 4142 9274
rect 4142 9222 4172 9274
rect 4196 9222 4206 9274
rect 4206 9222 4252 9274
rect 3956 9220 4012 9222
rect 4036 9220 4092 9222
rect 4116 9220 4172 9222
rect 4196 9220 4252 9222
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 938 5480 994 5536
rect 938 2796 940 2816
rect 940 2796 992 2816
rect 992 2796 994 2816
rect 938 2760 994 2796
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 4616 8730 4672 8732
rect 4696 8730 4752 8732
rect 4776 8730 4832 8732
rect 4856 8730 4912 8732
rect 4616 8678 4662 8730
rect 4662 8678 4672 8730
rect 4696 8678 4726 8730
rect 4726 8678 4738 8730
rect 4738 8678 4752 8730
rect 4776 8678 4790 8730
rect 4790 8678 4802 8730
rect 4802 8678 4832 8730
rect 4856 8678 4866 8730
rect 4866 8678 4912 8730
rect 4616 8676 4672 8678
rect 4696 8676 4752 8678
rect 4776 8676 4832 8678
rect 4856 8676 4912 8678
rect 5956 9274 6012 9276
rect 6036 9274 6092 9276
rect 6116 9274 6172 9276
rect 6196 9274 6252 9276
rect 5956 9222 6002 9274
rect 6002 9222 6012 9274
rect 6036 9222 6066 9274
rect 6066 9222 6078 9274
rect 6078 9222 6092 9274
rect 6116 9222 6130 9274
rect 6130 9222 6142 9274
rect 6142 9222 6172 9274
rect 6196 9222 6206 9274
rect 6206 9222 6252 9274
rect 5956 9220 6012 9222
rect 6036 9220 6092 9222
rect 6116 9220 6172 9222
rect 6196 9220 6252 9222
rect 3956 8186 4012 8188
rect 4036 8186 4092 8188
rect 4116 8186 4172 8188
rect 4196 8186 4252 8188
rect 3956 8134 4002 8186
rect 4002 8134 4012 8186
rect 4036 8134 4066 8186
rect 4066 8134 4078 8186
rect 4078 8134 4092 8186
rect 4116 8134 4130 8186
rect 4130 8134 4142 8186
rect 4142 8134 4172 8186
rect 4196 8134 4206 8186
rect 4206 8134 4252 8186
rect 3956 8132 4012 8134
rect 4036 8132 4092 8134
rect 4116 8132 4172 8134
rect 4196 8132 4252 8134
rect 4616 7642 4672 7644
rect 4696 7642 4752 7644
rect 4776 7642 4832 7644
rect 4856 7642 4912 7644
rect 4616 7590 4662 7642
rect 4662 7590 4672 7642
rect 4696 7590 4726 7642
rect 4726 7590 4738 7642
rect 4738 7590 4752 7642
rect 4776 7590 4790 7642
rect 4790 7590 4802 7642
rect 4802 7590 4832 7642
rect 4856 7590 4866 7642
rect 4866 7590 4912 7642
rect 4616 7588 4672 7590
rect 4696 7588 4752 7590
rect 4776 7588 4832 7590
rect 4856 7588 4912 7590
rect 3956 7098 4012 7100
rect 4036 7098 4092 7100
rect 4116 7098 4172 7100
rect 4196 7098 4252 7100
rect 3956 7046 4002 7098
rect 4002 7046 4012 7098
rect 4036 7046 4066 7098
rect 4066 7046 4078 7098
rect 4078 7046 4092 7098
rect 4116 7046 4130 7098
rect 4130 7046 4142 7098
rect 4142 7046 4172 7098
rect 4196 7046 4206 7098
rect 4206 7046 4252 7098
rect 3956 7044 4012 7046
rect 4036 7044 4092 7046
rect 4116 7044 4172 7046
rect 4196 7044 4252 7046
rect 4616 6554 4672 6556
rect 4696 6554 4752 6556
rect 4776 6554 4832 6556
rect 4856 6554 4912 6556
rect 4616 6502 4662 6554
rect 4662 6502 4672 6554
rect 4696 6502 4726 6554
rect 4726 6502 4738 6554
rect 4738 6502 4752 6554
rect 4776 6502 4790 6554
rect 4790 6502 4802 6554
rect 4802 6502 4832 6554
rect 4856 6502 4866 6554
rect 4866 6502 4912 6554
rect 4616 6500 4672 6502
rect 4696 6500 4752 6502
rect 4776 6500 4832 6502
rect 4856 6500 4912 6502
rect 3956 6010 4012 6012
rect 4036 6010 4092 6012
rect 4116 6010 4172 6012
rect 4196 6010 4252 6012
rect 3956 5958 4002 6010
rect 4002 5958 4012 6010
rect 4036 5958 4066 6010
rect 4066 5958 4078 6010
rect 4078 5958 4092 6010
rect 4116 5958 4130 6010
rect 4130 5958 4142 6010
rect 4142 5958 4172 6010
rect 4196 5958 4206 6010
rect 4206 5958 4252 6010
rect 3956 5956 4012 5958
rect 4036 5956 4092 5958
rect 4116 5956 4172 5958
rect 4196 5956 4252 5958
rect 4616 5466 4672 5468
rect 4696 5466 4752 5468
rect 4776 5466 4832 5468
rect 4856 5466 4912 5468
rect 4616 5414 4662 5466
rect 4662 5414 4672 5466
rect 4696 5414 4726 5466
rect 4726 5414 4738 5466
rect 4738 5414 4752 5466
rect 4776 5414 4790 5466
rect 4790 5414 4802 5466
rect 4802 5414 4832 5466
rect 4856 5414 4866 5466
rect 4866 5414 4912 5466
rect 4616 5412 4672 5414
rect 4696 5412 4752 5414
rect 4776 5412 4832 5414
rect 4856 5412 4912 5414
rect 3956 4922 4012 4924
rect 4036 4922 4092 4924
rect 4116 4922 4172 4924
rect 4196 4922 4252 4924
rect 3956 4870 4002 4922
rect 4002 4870 4012 4922
rect 4036 4870 4066 4922
rect 4066 4870 4078 4922
rect 4078 4870 4092 4922
rect 4116 4870 4130 4922
rect 4130 4870 4142 4922
rect 4142 4870 4172 4922
rect 4196 4870 4206 4922
rect 4206 4870 4252 4922
rect 3956 4868 4012 4870
rect 4036 4868 4092 4870
rect 4116 4868 4172 4870
rect 4196 4868 4252 4870
rect 3956 3834 4012 3836
rect 4036 3834 4092 3836
rect 4116 3834 4172 3836
rect 4196 3834 4252 3836
rect 3956 3782 4002 3834
rect 4002 3782 4012 3834
rect 4036 3782 4066 3834
rect 4066 3782 4078 3834
rect 4078 3782 4092 3834
rect 4116 3782 4130 3834
rect 4130 3782 4142 3834
rect 4142 3782 4172 3834
rect 4196 3782 4206 3834
rect 4206 3782 4252 3834
rect 3956 3780 4012 3782
rect 4036 3780 4092 3782
rect 4116 3780 4172 3782
rect 4196 3780 4252 3782
rect 4616 4378 4672 4380
rect 4696 4378 4752 4380
rect 4776 4378 4832 4380
rect 4856 4378 4912 4380
rect 4616 4326 4662 4378
rect 4662 4326 4672 4378
rect 4696 4326 4726 4378
rect 4726 4326 4738 4378
rect 4738 4326 4752 4378
rect 4776 4326 4790 4378
rect 4790 4326 4802 4378
rect 4802 4326 4832 4378
rect 4856 4326 4866 4378
rect 4866 4326 4912 4378
rect 4616 4324 4672 4326
rect 4696 4324 4752 4326
rect 4776 4324 4832 4326
rect 4856 4324 4912 4326
rect 4616 3290 4672 3292
rect 4696 3290 4752 3292
rect 4776 3290 4832 3292
rect 4856 3290 4912 3292
rect 4616 3238 4662 3290
rect 4662 3238 4672 3290
rect 4696 3238 4726 3290
rect 4726 3238 4738 3290
rect 4738 3238 4752 3290
rect 4776 3238 4790 3290
rect 4790 3238 4802 3290
rect 4802 3238 4832 3290
rect 4856 3238 4866 3290
rect 4866 3238 4912 3290
rect 4616 3236 4672 3238
rect 4696 3236 4752 3238
rect 4776 3236 4832 3238
rect 4856 3236 4912 3238
rect 6616 8730 6672 8732
rect 6696 8730 6752 8732
rect 6776 8730 6832 8732
rect 6856 8730 6912 8732
rect 6616 8678 6662 8730
rect 6662 8678 6672 8730
rect 6696 8678 6726 8730
rect 6726 8678 6738 8730
rect 6738 8678 6752 8730
rect 6776 8678 6790 8730
rect 6790 8678 6802 8730
rect 6802 8678 6832 8730
rect 6856 8678 6866 8730
rect 6866 8678 6912 8730
rect 6616 8676 6672 8678
rect 6696 8676 6752 8678
rect 6776 8676 6832 8678
rect 6856 8676 6912 8678
rect 5956 8186 6012 8188
rect 6036 8186 6092 8188
rect 6116 8186 6172 8188
rect 6196 8186 6252 8188
rect 5956 8134 6002 8186
rect 6002 8134 6012 8186
rect 6036 8134 6066 8186
rect 6066 8134 6078 8186
rect 6078 8134 6092 8186
rect 6116 8134 6130 8186
rect 6130 8134 6142 8186
rect 6142 8134 6172 8186
rect 6196 8134 6206 8186
rect 6206 8134 6252 8186
rect 5956 8132 6012 8134
rect 6036 8132 6092 8134
rect 6116 8132 6172 8134
rect 6196 8132 6252 8134
rect 8942 9580 8998 9616
rect 8942 9560 8944 9580
rect 8944 9560 8996 9580
rect 8996 9560 8998 9580
rect 6616 7642 6672 7644
rect 6696 7642 6752 7644
rect 6776 7642 6832 7644
rect 6856 7642 6912 7644
rect 6616 7590 6662 7642
rect 6662 7590 6672 7642
rect 6696 7590 6726 7642
rect 6726 7590 6738 7642
rect 6738 7590 6752 7642
rect 6776 7590 6790 7642
rect 6790 7590 6802 7642
rect 6802 7590 6832 7642
rect 6856 7590 6866 7642
rect 6866 7590 6912 7642
rect 6616 7588 6672 7590
rect 6696 7588 6752 7590
rect 6776 7588 6832 7590
rect 6856 7588 6912 7590
rect 5956 7098 6012 7100
rect 6036 7098 6092 7100
rect 6116 7098 6172 7100
rect 6196 7098 6252 7100
rect 5956 7046 6002 7098
rect 6002 7046 6012 7098
rect 6036 7046 6066 7098
rect 6066 7046 6078 7098
rect 6078 7046 6092 7098
rect 6116 7046 6130 7098
rect 6130 7046 6142 7098
rect 6142 7046 6172 7098
rect 6196 7046 6206 7098
rect 6206 7046 6252 7098
rect 5956 7044 6012 7046
rect 6036 7044 6092 7046
rect 6116 7044 6172 7046
rect 6196 7044 6252 7046
rect 5956 6010 6012 6012
rect 6036 6010 6092 6012
rect 6116 6010 6172 6012
rect 6196 6010 6252 6012
rect 5956 5958 6002 6010
rect 6002 5958 6012 6010
rect 6036 5958 6066 6010
rect 6066 5958 6078 6010
rect 6078 5958 6092 6010
rect 6116 5958 6130 6010
rect 6130 5958 6142 6010
rect 6142 5958 6172 6010
rect 6196 5958 6206 6010
rect 6206 5958 6252 6010
rect 5956 5956 6012 5958
rect 6036 5956 6092 5958
rect 6116 5956 6172 5958
rect 6196 5956 6252 5958
rect 5956 4922 6012 4924
rect 6036 4922 6092 4924
rect 6116 4922 6172 4924
rect 6196 4922 6252 4924
rect 5956 4870 6002 4922
rect 6002 4870 6012 4922
rect 6036 4870 6066 4922
rect 6066 4870 6078 4922
rect 6078 4870 6092 4922
rect 6116 4870 6130 4922
rect 6130 4870 6142 4922
rect 6142 4870 6172 4922
rect 6196 4870 6206 4922
rect 6206 4870 6252 4922
rect 5956 4868 6012 4870
rect 6036 4868 6092 4870
rect 6116 4868 6172 4870
rect 6196 4868 6252 4870
rect 5956 3834 6012 3836
rect 6036 3834 6092 3836
rect 6116 3834 6172 3836
rect 6196 3834 6252 3836
rect 5956 3782 6002 3834
rect 6002 3782 6012 3834
rect 6036 3782 6066 3834
rect 6066 3782 6078 3834
rect 6078 3782 6092 3834
rect 6116 3782 6130 3834
rect 6130 3782 6142 3834
rect 6142 3782 6172 3834
rect 6196 3782 6206 3834
rect 6206 3782 6252 3834
rect 5956 3780 6012 3782
rect 6036 3780 6092 3782
rect 6116 3780 6172 3782
rect 6196 3780 6252 3782
rect 6616 6554 6672 6556
rect 6696 6554 6752 6556
rect 6776 6554 6832 6556
rect 6856 6554 6912 6556
rect 6616 6502 6662 6554
rect 6662 6502 6672 6554
rect 6696 6502 6726 6554
rect 6726 6502 6738 6554
rect 6738 6502 6752 6554
rect 6776 6502 6790 6554
rect 6790 6502 6802 6554
rect 6802 6502 6832 6554
rect 6856 6502 6866 6554
rect 6866 6502 6912 6554
rect 6616 6500 6672 6502
rect 6696 6500 6752 6502
rect 6776 6500 6832 6502
rect 6856 6500 6912 6502
rect 7956 9274 8012 9276
rect 8036 9274 8092 9276
rect 8116 9274 8172 9276
rect 8196 9274 8252 9276
rect 7956 9222 8002 9274
rect 8002 9222 8012 9274
rect 8036 9222 8066 9274
rect 8066 9222 8078 9274
rect 8078 9222 8092 9274
rect 8116 9222 8130 9274
rect 8130 9222 8142 9274
rect 8142 9222 8172 9274
rect 8196 9222 8206 9274
rect 8206 9222 8252 9274
rect 7956 9220 8012 9222
rect 8036 9220 8092 9222
rect 8116 9220 8172 9222
rect 8196 9220 8252 9222
rect 8616 8730 8672 8732
rect 8696 8730 8752 8732
rect 8776 8730 8832 8732
rect 8856 8730 8912 8732
rect 8616 8678 8662 8730
rect 8662 8678 8672 8730
rect 8696 8678 8726 8730
rect 8726 8678 8738 8730
rect 8738 8678 8752 8730
rect 8776 8678 8790 8730
rect 8790 8678 8802 8730
rect 8802 8678 8832 8730
rect 8856 8678 8866 8730
rect 8866 8678 8912 8730
rect 8616 8676 8672 8678
rect 8696 8676 8752 8678
rect 8776 8676 8832 8678
rect 8856 8676 8912 8678
rect 7956 8186 8012 8188
rect 8036 8186 8092 8188
rect 8116 8186 8172 8188
rect 8196 8186 8252 8188
rect 7956 8134 8002 8186
rect 8002 8134 8012 8186
rect 8036 8134 8066 8186
rect 8066 8134 8078 8186
rect 8078 8134 8092 8186
rect 8116 8134 8130 8186
rect 8130 8134 8142 8186
rect 8142 8134 8172 8186
rect 8196 8134 8206 8186
rect 8206 8134 8252 8186
rect 7956 8132 8012 8134
rect 8036 8132 8092 8134
rect 8116 8132 8172 8134
rect 8196 8132 8252 8134
rect 8616 7642 8672 7644
rect 8696 7642 8752 7644
rect 8776 7642 8832 7644
rect 8856 7642 8912 7644
rect 8616 7590 8662 7642
rect 8662 7590 8672 7642
rect 8696 7590 8726 7642
rect 8726 7590 8738 7642
rect 8738 7590 8752 7642
rect 8776 7590 8790 7642
rect 8790 7590 8802 7642
rect 8802 7590 8832 7642
rect 8856 7590 8866 7642
rect 8866 7590 8912 7642
rect 8616 7588 8672 7590
rect 8696 7588 8752 7590
rect 8776 7588 8832 7590
rect 8856 7588 8912 7590
rect 7956 7098 8012 7100
rect 8036 7098 8092 7100
rect 8116 7098 8172 7100
rect 8196 7098 8252 7100
rect 7956 7046 8002 7098
rect 8002 7046 8012 7098
rect 8036 7046 8066 7098
rect 8066 7046 8078 7098
rect 8078 7046 8092 7098
rect 8116 7046 8130 7098
rect 8130 7046 8142 7098
rect 8142 7046 8172 7098
rect 8196 7046 8206 7098
rect 8206 7046 8252 7098
rect 7956 7044 8012 7046
rect 8036 7044 8092 7046
rect 8116 7044 8172 7046
rect 8196 7044 8252 7046
rect 9218 6840 9274 6896
rect 8616 6554 8672 6556
rect 8696 6554 8752 6556
rect 8776 6554 8832 6556
rect 8856 6554 8912 6556
rect 8616 6502 8662 6554
rect 8662 6502 8672 6554
rect 8696 6502 8726 6554
rect 8726 6502 8738 6554
rect 8738 6502 8752 6554
rect 8776 6502 8790 6554
rect 8790 6502 8802 6554
rect 8802 6502 8832 6554
rect 8856 6502 8866 6554
rect 8866 6502 8912 6554
rect 8616 6500 8672 6502
rect 8696 6500 8752 6502
rect 8776 6500 8832 6502
rect 8856 6500 8912 6502
rect 7956 6010 8012 6012
rect 8036 6010 8092 6012
rect 8116 6010 8172 6012
rect 8196 6010 8252 6012
rect 7956 5958 8002 6010
rect 8002 5958 8012 6010
rect 8036 5958 8066 6010
rect 8066 5958 8078 6010
rect 8078 5958 8092 6010
rect 8116 5958 8130 6010
rect 8130 5958 8142 6010
rect 8142 5958 8172 6010
rect 8196 5958 8206 6010
rect 8206 5958 8252 6010
rect 7956 5956 8012 5958
rect 8036 5956 8092 5958
rect 8116 5956 8172 5958
rect 8196 5956 8252 5958
rect 6616 5466 6672 5468
rect 6696 5466 6752 5468
rect 6776 5466 6832 5468
rect 6856 5466 6912 5468
rect 6616 5414 6662 5466
rect 6662 5414 6672 5466
rect 6696 5414 6726 5466
rect 6726 5414 6738 5466
rect 6738 5414 6752 5466
rect 6776 5414 6790 5466
rect 6790 5414 6802 5466
rect 6802 5414 6832 5466
rect 6856 5414 6866 5466
rect 6866 5414 6912 5466
rect 6616 5412 6672 5414
rect 6696 5412 6752 5414
rect 6776 5412 6832 5414
rect 6856 5412 6912 5414
rect 6616 4378 6672 4380
rect 6696 4378 6752 4380
rect 6776 4378 6832 4380
rect 6856 4378 6912 4380
rect 6616 4326 6662 4378
rect 6662 4326 6672 4378
rect 6696 4326 6726 4378
rect 6726 4326 6738 4378
rect 6738 4326 6752 4378
rect 6776 4326 6790 4378
rect 6790 4326 6802 4378
rect 6802 4326 6832 4378
rect 6856 4326 6866 4378
rect 6866 4326 6912 4378
rect 6616 4324 6672 4326
rect 6696 4324 6752 4326
rect 6776 4324 6832 4326
rect 6856 4324 6912 4326
rect 7956 4922 8012 4924
rect 8036 4922 8092 4924
rect 8116 4922 8172 4924
rect 8196 4922 8252 4924
rect 7956 4870 8002 4922
rect 8002 4870 8012 4922
rect 8036 4870 8066 4922
rect 8066 4870 8078 4922
rect 8078 4870 8092 4922
rect 8116 4870 8130 4922
rect 8130 4870 8142 4922
rect 8142 4870 8172 4922
rect 8196 4870 8206 4922
rect 8206 4870 8252 4922
rect 7956 4868 8012 4870
rect 8036 4868 8092 4870
rect 8116 4868 8172 4870
rect 8196 4868 8252 4870
rect 6616 3290 6672 3292
rect 6696 3290 6752 3292
rect 6776 3290 6832 3292
rect 6856 3290 6912 3292
rect 6616 3238 6662 3290
rect 6662 3238 6672 3290
rect 6696 3238 6726 3290
rect 6726 3238 6738 3290
rect 6738 3238 6752 3290
rect 6776 3238 6790 3290
rect 6790 3238 6802 3290
rect 6802 3238 6832 3290
rect 6856 3238 6866 3290
rect 6866 3238 6912 3290
rect 6616 3236 6672 3238
rect 6696 3236 6752 3238
rect 6776 3236 6832 3238
rect 6856 3236 6912 3238
rect 7956 3834 8012 3836
rect 8036 3834 8092 3836
rect 8116 3834 8172 3836
rect 8196 3834 8252 3836
rect 7956 3782 8002 3834
rect 8002 3782 8012 3834
rect 8036 3782 8066 3834
rect 8066 3782 8078 3834
rect 8078 3782 8092 3834
rect 8116 3782 8130 3834
rect 8130 3782 8142 3834
rect 8142 3782 8172 3834
rect 8196 3782 8206 3834
rect 8206 3782 8252 3834
rect 7956 3780 8012 3782
rect 8036 3780 8092 3782
rect 8116 3780 8172 3782
rect 8196 3780 8252 3782
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 3956 2746 4012 2748
rect 4036 2746 4092 2748
rect 4116 2746 4172 2748
rect 4196 2746 4252 2748
rect 3956 2694 4002 2746
rect 4002 2694 4012 2746
rect 4036 2694 4066 2746
rect 4066 2694 4078 2746
rect 4078 2694 4092 2746
rect 4116 2694 4130 2746
rect 4130 2694 4142 2746
rect 4142 2694 4172 2746
rect 4196 2694 4206 2746
rect 4206 2694 4252 2746
rect 3956 2692 4012 2694
rect 4036 2692 4092 2694
rect 4116 2692 4172 2694
rect 4196 2692 4252 2694
rect 5956 2746 6012 2748
rect 6036 2746 6092 2748
rect 6116 2746 6172 2748
rect 6196 2746 6252 2748
rect 5956 2694 6002 2746
rect 6002 2694 6012 2746
rect 6036 2694 6066 2746
rect 6066 2694 6078 2746
rect 6078 2694 6092 2746
rect 6116 2694 6130 2746
rect 6130 2694 6142 2746
rect 6142 2694 6172 2746
rect 6196 2694 6206 2746
rect 6206 2694 6252 2746
rect 5956 2692 6012 2694
rect 6036 2692 6092 2694
rect 6116 2692 6172 2694
rect 6196 2692 6252 2694
rect 7956 2746 8012 2748
rect 8036 2746 8092 2748
rect 8116 2746 8172 2748
rect 8196 2746 8252 2748
rect 7956 2694 8002 2746
rect 8002 2694 8012 2746
rect 8036 2694 8066 2746
rect 8066 2694 8078 2746
rect 8078 2694 8092 2746
rect 8116 2694 8130 2746
rect 8130 2694 8142 2746
rect 8142 2694 8172 2746
rect 8196 2694 8206 2746
rect 8206 2694 8252 2746
rect 7956 2692 8012 2694
rect 8036 2692 8092 2694
rect 8116 2692 8172 2694
rect 8196 2692 8252 2694
rect 8616 5466 8672 5468
rect 8696 5466 8752 5468
rect 8776 5466 8832 5468
rect 8856 5466 8912 5468
rect 8616 5414 8662 5466
rect 8662 5414 8672 5466
rect 8696 5414 8726 5466
rect 8726 5414 8738 5466
rect 8738 5414 8752 5466
rect 8776 5414 8790 5466
rect 8790 5414 8802 5466
rect 8802 5414 8832 5466
rect 8856 5414 8866 5466
rect 8866 5414 8912 5466
rect 8616 5412 8672 5414
rect 8696 5412 8752 5414
rect 8776 5412 8832 5414
rect 8856 5412 8912 5414
rect 8616 4378 8672 4380
rect 8696 4378 8752 4380
rect 8776 4378 8832 4380
rect 8856 4378 8912 4380
rect 8616 4326 8662 4378
rect 8662 4326 8672 4378
rect 8696 4326 8726 4378
rect 8726 4326 8738 4378
rect 8738 4326 8752 4378
rect 8776 4326 8790 4378
rect 8790 4326 8802 4378
rect 8802 4326 8832 4378
rect 8856 4326 8866 4378
rect 8866 4326 8912 4378
rect 8616 4324 8672 4326
rect 8696 4324 8752 4326
rect 8776 4324 8832 4326
rect 8856 4324 8912 4326
rect 9218 3476 9220 3496
rect 9220 3476 9272 3496
rect 9272 3476 9274 3496
rect 9218 3440 9274 3476
rect 8616 3290 8672 3292
rect 8696 3290 8752 3292
rect 8776 3290 8832 3292
rect 8856 3290 8912 3292
rect 8616 3238 8662 3290
rect 8662 3238 8672 3290
rect 8696 3238 8726 3290
rect 8726 3238 8738 3290
rect 8738 3238 8752 3290
rect 8776 3238 8790 3290
rect 8790 3238 8802 3290
rect 8802 3238 8832 3290
rect 8856 3238 8866 3290
rect 8866 3238 8912 3290
rect 8616 3236 8672 3238
rect 8696 3236 8752 3238
rect 8776 3236 8832 3238
rect 8856 3236 8912 3238
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 4616 2202 4672 2204
rect 4696 2202 4752 2204
rect 4776 2202 4832 2204
rect 4856 2202 4912 2204
rect 4616 2150 4662 2202
rect 4662 2150 4672 2202
rect 4696 2150 4726 2202
rect 4726 2150 4738 2202
rect 4738 2150 4752 2202
rect 4776 2150 4790 2202
rect 4790 2150 4802 2202
rect 4802 2150 4832 2202
rect 4856 2150 4866 2202
rect 4866 2150 4912 2202
rect 4616 2148 4672 2150
rect 4696 2148 4752 2150
rect 4776 2148 4832 2150
rect 4856 2148 4912 2150
rect 6616 2202 6672 2204
rect 6696 2202 6752 2204
rect 6776 2202 6832 2204
rect 6856 2202 6912 2204
rect 6616 2150 6662 2202
rect 6662 2150 6672 2202
rect 6696 2150 6726 2202
rect 6726 2150 6738 2202
rect 6738 2150 6752 2202
rect 6776 2150 6790 2202
rect 6790 2150 6802 2202
rect 6802 2150 6832 2202
rect 6856 2150 6866 2202
rect 6866 2150 6912 2202
rect 6616 2148 6672 2150
rect 6696 2148 6752 2150
rect 6776 2148 6832 2150
rect 6856 2148 6912 2150
rect 8616 2202 8672 2204
rect 8696 2202 8752 2204
rect 8776 2202 8832 2204
rect 8856 2202 8912 2204
rect 8616 2150 8662 2202
rect 8662 2150 8672 2202
rect 8696 2150 8726 2202
rect 8726 2150 8738 2202
rect 8738 2150 8752 2202
rect 8776 2150 8790 2202
rect 8790 2150 8802 2202
rect 8802 2150 8832 2202
rect 8856 2150 8866 2202
rect 8866 2150 8912 2202
rect 8616 2148 8672 2150
rect 8696 2148 8752 2150
rect 8776 2148 8832 2150
rect 8856 2148 8912 2150
rect 9034 720 9090 776
<< metal3 >>
rect 0 11658 800 11688
rect 0 11598 1042 11658
rect 0 11568 800 11598
rect 982 11386 1042 11598
rect 1853 11386 1919 11389
rect 982 11384 1919 11386
rect 982 11328 1858 11384
rect 1914 11328 1919 11384
rect 982 11326 1919 11328
rect 1853 11323 1919 11326
rect 2606 9824 2922 9825
rect 2606 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2922 9824
rect 2606 9759 2922 9760
rect 4606 9824 4922 9825
rect 4606 9760 4612 9824
rect 4676 9760 4692 9824
rect 4756 9760 4772 9824
rect 4836 9760 4852 9824
rect 4916 9760 4922 9824
rect 4606 9759 4922 9760
rect 6606 9824 6922 9825
rect 6606 9760 6612 9824
rect 6676 9760 6692 9824
rect 6756 9760 6772 9824
rect 6836 9760 6852 9824
rect 6916 9760 6922 9824
rect 6606 9759 6922 9760
rect 8606 9824 8922 9825
rect 8606 9760 8612 9824
rect 8676 9760 8692 9824
rect 8756 9760 8772 9824
rect 8836 9760 8852 9824
rect 8916 9760 8922 9824
rect 8606 9759 8922 9760
rect 8937 9618 9003 9621
rect 9474 9618 10274 9648
rect 8937 9616 10274 9618
rect 8937 9560 8942 9616
rect 8998 9560 10274 9616
rect 8937 9558 10274 9560
rect 8937 9555 9003 9558
rect 9474 9528 10274 9558
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 3946 9280 4262 9281
rect 3946 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4112 9280
rect 4176 9216 4192 9280
rect 4256 9216 4262 9280
rect 3946 9215 4262 9216
rect 5946 9280 6262 9281
rect 5946 9216 5952 9280
rect 6016 9216 6032 9280
rect 6096 9216 6112 9280
rect 6176 9216 6192 9280
rect 6256 9216 6262 9280
rect 5946 9215 6262 9216
rect 7946 9280 8262 9281
rect 7946 9216 7952 9280
rect 8016 9216 8032 9280
rect 8096 9216 8112 9280
rect 8176 9216 8192 9280
rect 8256 9216 8262 9280
rect 7946 9215 8262 9216
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 4606 8736 4922 8737
rect 4606 8672 4612 8736
rect 4676 8672 4692 8736
rect 4756 8672 4772 8736
rect 4836 8672 4852 8736
rect 4916 8672 4922 8736
rect 4606 8671 4922 8672
rect 6606 8736 6922 8737
rect 6606 8672 6612 8736
rect 6676 8672 6692 8736
rect 6756 8672 6772 8736
rect 6836 8672 6852 8736
rect 6916 8672 6922 8736
rect 6606 8671 6922 8672
rect 8606 8736 8922 8737
rect 8606 8672 8612 8736
rect 8676 8672 8692 8736
rect 8756 8672 8772 8736
rect 8836 8672 8852 8736
rect 8916 8672 8922 8736
rect 8606 8671 8922 8672
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 3946 8192 4262 8193
rect 3946 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4112 8192
rect 4176 8128 4192 8192
rect 4256 8128 4262 8192
rect 3946 8127 4262 8128
rect 5946 8192 6262 8193
rect 5946 8128 5952 8192
rect 6016 8128 6032 8192
rect 6096 8128 6112 8192
rect 6176 8128 6192 8192
rect 6256 8128 6262 8192
rect 5946 8127 6262 8128
rect 7946 8192 8262 8193
rect 7946 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8262 8192
rect 7946 8127 8262 8128
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 2606 7583 2922 7584
rect 4606 7648 4922 7649
rect 4606 7584 4612 7648
rect 4676 7584 4692 7648
rect 4756 7584 4772 7648
rect 4836 7584 4852 7648
rect 4916 7584 4922 7648
rect 4606 7583 4922 7584
rect 6606 7648 6922 7649
rect 6606 7584 6612 7648
rect 6676 7584 6692 7648
rect 6756 7584 6772 7648
rect 6836 7584 6852 7648
rect 6916 7584 6922 7648
rect 6606 7583 6922 7584
rect 8606 7648 8922 7649
rect 8606 7584 8612 7648
rect 8676 7584 8692 7648
rect 8756 7584 8772 7648
rect 8836 7584 8852 7648
rect 8916 7584 8922 7648
rect 8606 7583 8922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 3946 7104 4262 7105
rect 3946 7040 3952 7104
rect 4016 7040 4032 7104
rect 4096 7040 4112 7104
rect 4176 7040 4192 7104
rect 4256 7040 4262 7104
rect 3946 7039 4262 7040
rect 5946 7104 6262 7105
rect 5946 7040 5952 7104
rect 6016 7040 6032 7104
rect 6096 7040 6112 7104
rect 6176 7040 6192 7104
rect 6256 7040 6262 7104
rect 5946 7039 6262 7040
rect 7946 7104 8262 7105
rect 7946 7040 7952 7104
rect 8016 7040 8032 7104
rect 8096 7040 8112 7104
rect 8176 7040 8192 7104
rect 8256 7040 8262 7104
rect 7946 7039 8262 7040
rect 9213 6898 9279 6901
rect 9474 6898 10274 6928
rect 9213 6896 10274 6898
rect 9213 6840 9218 6896
rect 9274 6840 10274 6896
rect 9213 6838 10274 6840
rect 9213 6835 9279 6838
rect 9474 6808 10274 6838
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 4606 6560 4922 6561
rect 4606 6496 4612 6560
rect 4676 6496 4692 6560
rect 4756 6496 4772 6560
rect 4836 6496 4852 6560
rect 4916 6496 4922 6560
rect 4606 6495 4922 6496
rect 6606 6560 6922 6561
rect 6606 6496 6612 6560
rect 6676 6496 6692 6560
rect 6756 6496 6772 6560
rect 6836 6496 6852 6560
rect 6916 6496 6922 6560
rect 6606 6495 6922 6496
rect 8606 6560 8922 6561
rect 8606 6496 8612 6560
rect 8676 6496 8692 6560
rect 8756 6496 8772 6560
rect 8836 6496 8852 6560
rect 8916 6496 8922 6560
rect 8606 6495 8922 6496
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 3946 6016 4262 6017
rect 3946 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4112 6016
rect 4176 5952 4192 6016
rect 4256 5952 4262 6016
rect 3946 5951 4262 5952
rect 5946 6016 6262 6017
rect 5946 5952 5952 6016
rect 6016 5952 6032 6016
rect 6096 5952 6112 6016
rect 6176 5952 6192 6016
rect 6256 5952 6262 6016
rect 5946 5951 6262 5952
rect 7946 6016 8262 6017
rect 7946 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8262 6016
rect 7946 5951 8262 5952
rect 0 5538 800 5568
rect 933 5538 999 5541
rect 0 5536 999 5538
rect 0 5480 938 5536
rect 994 5480 999 5536
rect 0 5478 999 5480
rect 0 5448 800 5478
rect 933 5475 999 5478
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 4606 5472 4922 5473
rect 4606 5408 4612 5472
rect 4676 5408 4692 5472
rect 4756 5408 4772 5472
rect 4836 5408 4852 5472
rect 4916 5408 4922 5472
rect 4606 5407 4922 5408
rect 6606 5472 6922 5473
rect 6606 5408 6612 5472
rect 6676 5408 6692 5472
rect 6756 5408 6772 5472
rect 6836 5408 6852 5472
rect 6916 5408 6922 5472
rect 6606 5407 6922 5408
rect 8606 5472 8922 5473
rect 8606 5408 8612 5472
rect 8676 5408 8692 5472
rect 8756 5408 8772 5472
rect 8836 5408 8852 5472
rect 8916 5408 8922 5472
rect 8606 5407 8922 5408
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 1946 4863 2262 4864
rect 3946 4928 4262 4929
rect 3946 4864 3952 4928
rect 4016 4864 4032 4928
rect 4096 4864 4112 4928
rect 4176 4864 4192 4928
rect 4256 4864 4262 4928
rect 3946 4863 4262 4864
rect 5946 4928 6262 4929
rect 5946 4864 5952 4928
rect 6016 4864 6032 4928
rect 6096 4864 6112 4928
rect 6176 4864 6192 4928
rect 6256 4864 6262 4928
rect 5946 4863 6262 4864
rect 7946 4928 8262 4929
rect 7946 4864 7952 4928
rect 8016 4864 8032 4928
rect 8096 4864 8112 4928
rect 8176 4864 8192 4928
rect 8256 4864 8262 4928
rect 7946 4863 8262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 4606 4384 4922 4385
rect 4606 4320 4612 4384
rect 4676 4320 4692 4384
rect 4756 4320 4772 4384
rect 4836 4320 4852 4384
rect 4916 4320 4922 4384
rect 4606 4319 4922 4320
rect 6606 4384 6922 4385
rect 6606 4320 6612 4384
rect 6676 4320 6692 4384
rect 6756 4320 6772 4384
rect 6836 4320 6852 4384
rect 6916 4320 6922 4384
rect 6606 4319 6922 4320
rect 8606 4384 8922 4385
rect 8606 4320 8612 4384
rect 8676 4320 8692 4384
rect 8756 4320 8772 4384
rect 8836 4320 8852 4384
rect 8916 4320 8922 4384
rect 8606 4319 8922 4320
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 3946 3840 4262 3841
rect 3946 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4112 3840
rect 4176 3776 4192 3840
rect 4256 3776 4262 3840
rect 3946 3775 4262 3776
rect 5946 3840 6262 3841
rect 5946 3776 5952 3840
rect 6016 3776 6032 3840
rect 6096 3776 6112 3840
rect 6176 3776 6192 3840
rect 6256 3776 6262 3840
rect 5946 3775 6262 3776
rect 7946 3840 8262 3841
rect 7946 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8262 3840
rect 7946 3775 8262 3776
rect 9213 3498 9279 3501
rect 9474 3498 10274 3528
rect 9213 3496 10274 3498
rect 9213 3440 9218 3496
rect 9274 3440 10274 3496
rect 9213 3438 10274 3440
rect 9213 3435 9279 3438
rect 9474 3408 10274 3438
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 4606 3296 4922 3297
rect 4606 3232 4612 3296
rect 4676 3232 4692 3296
rect 4756 3232 4772 3296
rect 4836 3232 4852 3296
rect 4916 3232 4922 3296
rect 4606 3231 4922 3232
rect 6606 3296 6922 3297
rect 6606 3232 6612 3296
rect 6676 3232 6692 3296
rect 6756 3232 6772 3296
rect 6836 3232 6852 3296
rect 6916 3232 6922 3296
rect 6606 3231 6922 3232
rect 8606 3296 8922 3297
rect 8606 3232 8612 3296
rect 8676 3232 8692 3296
rect 8756 3232 8772 3296
rect 8836 3232 8852 3296
rect 8916 3232 8922 3296
rect 8606 3231 8922 3232
rect 0 2818 800 2848
rect 933 2818 999 2821
rect 0 2816 999 2818
rect 0 2760 938 2816
rect 994 2760 999 2816
rect 0 2758 999 2760
rect 0 2728 800 2758
rect 933 2755 999 2758
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 3946 2752 4262 2753
rect 3946 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4112 2752
rect 4176 2688 4192 2752
rect 4256 2688 4262 2752
rect 3946 2687 4262 2688
rect 5946 2752 6262 2753
rect 5946 2688 5952 2752
rect 6016 2688 6032 2752
rect 6096 2688 6112 2752
rect 6176 2688 6192 2752
rect 6256 2688 6262 2752
rect 5946 2687 6262 2688
rect 7946 2752 8262 2753
rect 7946 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8262 2752
rect 7946 2687 8262 2688
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 2606 2143 2922 2144
rect 4606 2208 4922 2209
rect 4606 2144 4612 2208
rect 4676 2144 4692 2208
rect 4756 2144 4772 2208
rect 4836 2144 4852 2208
rect 4916 2144 4922 2208
rect 4606 2143 4922 2144
rect 6606 2208 6922 2209
rect 6606 2144 6612 2208
rect 6676 2144 6692 2208
rect 6756 2144 6772 2208
rect 6836 2144 6852 2208
rect 6916 2144 6922 2208
rect 6606 2143 6922 2144
rect 8606 2208 8922 2209
rect 8606 2144 8612 2208
rect 8676 2144 8692 2208
rect 8756 2144 8772 2208
rect 8836 2144 8852 2208
rect 8916 2144 8922 2208
rect 8606 2143 8922 2144
rect 9029 778 9095 781
rect 9474 778 10274 808
rect 9029 776 10274 778
rect 9029 720 9034 776
rect 9090 720 10274 776
rect 9029 718 10274 720
rect 9029 715 9095 718
rect 9474 688 10274 718
<< via3 >>
rect 2612 9820 2676 9824
rect 2612 9764 2616 9820
rect 2616 9764 2672 9820
rect 2672 9764 2676 9820
rect 2612 9760 2676 9764
rect 2692 9820 2756 9824
rect 2692 9764 2696 9820
rect 2696 9764 2752 9820
rect 2752 9764 2756 9820
rect 2692 9760 2756 9764
rect 2772 9820 2836 9824
rect 2772 9764 2776 9820
rect 2776 9764 2832 9820
rect 2832 9764 2836 9820
rect 2772 9760 2836 9764
rect 2852 9820 2916 9824
rect 2852 9764 2856 9820
rect 2856 9764 2912 9820
rect 2912 9764 2916 9820
rect 2852 9760 2916 9764
rect 4612 9820 4676 9824
rect 4612 9764 4616 9820
rect 4616 9764 4672 9820
rect 4672 9764 4676 9820
rect 4612 9760 4676 9764
rect 4692 9820 4756 9824
rect 4692 9764 4696 9820
rect 4696 9764 4752 9820
rect 4752 9764 4756 9820
rect 4692 9760 4756 9764
rect 4772 9820 4836 9824
rect 4772 9764 4776 9820
rect 4776 9764 4832 9820
rect 4832 9764 4836 9820
rect 4772 9760 4836 9764
rect 4852 9820 4916 9824
rect 4852 9764 4856 9820
rect 4856 9764 4912 9820
rect 4912 9764 4916 9820
rect 4852 9760 4916 9764
rect 6612 9820 6676 9824
rect 6612 9764 6616 9820
rect 6616 9764 6672 9820
rect 6672 9764 6676 9820
rect 6612 9760 6676 9764
rect 6692 9820 6756 9824
rect 6692 9764 6696 9820
rect 6696 9764 6752 9820
rect 6752 9764 6756 9820
rect 6692 9760 6756 9764
rect 6772 9820 6836 9824
rect 6772 9764 6776 9820
rect 6776 9764 6832 9820
rect 6832 9764 6836 9820
rect 6772 9760 6836 9764
rect 6852 9820 6916 9824
rect 6852 9764 6856 9820
rect 6856 9764 6912 9820
rect 6912 9764 6916 9820
rect 6852 9760 6916 9764
rect 8612 9820 8676 9824
rect 8612 9764 8616 9820
rect 8616 9764 8672 9820
rect 8672 9764 8676 9820
rect 8612 9760 8676 9764
rect 8692 9820 8756 9824
rect 8692 9764 8696 9820
rect 8696 9764 8752 9820
rect 8752 9764 8756 9820
rect 8692 9760 8756 9764
rect 8772 9820 8836 9824
rect 8772 9764 8776 9820
rect 8776 9764 8832 9820
rect 8832 9764 8836 9820
rect 8772 9760 8836 9764
rect 8852 9820 8916 9824
rect 8852 9764 8856 9820
rect 8856 9764 8912 9820
rect 8912 9764 8916 9820
rect 8852 9760 8916 9764
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 3952 9276 4016 9280
rect 3952 9220 3956 9276
rect 3956 9220 4012 9276
rect 4012 9220 4016 9276
rect 3952 9216 4016 9220
rect 4032 9276 4096 9280
rect 4032 9220 4036 9276
rect 4036 9220 4092 9276
rect 4092 9220 4096 9276
rect 4032 9216 4096 9220
rect 4112 9276 4176 9280
rect 4112 9220 4116 9276
rect 4116 9220 4172 9276
rect 4172 9220 4176 9276
rect 4112 9216 4176 9220
rect 4192 9276 4256 9280
rect 4192 9220 4196 9276
rect 4196 9220 4252 9276
rect 4252 9220 4256 9276
rect 4192 9216 4256 9220
rect 5952 9276 6016 9280
rect 5952 9220 5956 9276
rect 5956 9220 6012 9276
rect 6012 9220 6016 9276
rect 5952 9216 6016 9220
rect 6032 9276 6096 9280
rect 6032 9220 6036 9276
rect 6036 9220 6092 9276
rect 6092 9220 6096 9276
rect 6032 9216 6096 9220
rect 6112 9276 6176 9280
rect 6112 9220 6116 9276
rect 6116 9220 6172 9276
rect 6172 9220 6176 9276
rect 6112 9216 6176 9220
rect 6192 9276 6256 9280
rect 6192 9220 6196 9276
rect 6196 9220 6252 9276
rect 6252 9220 6256 9276
rect 6192 9216 6256 9220
rect 7952 9276 8016 9280
rect 7952 9220 7956 9276
rect 7956 9220 8012 9276
rect 8012 9220 8016 9276
rect 7952 9216 8016 9220
rect 8032 9276 8096 9280
rect 8032 9220 8036 9276
rect 8036 9220 8092 9276
rect 8092 9220 8096 9276
rect 8032 9216 8096 9220
rect 8112 9276 8176 9280
rect 8112 9220 8116 9276
rect 8116 9220 8172 9276
rect 8172 9220 8176 9276
rect 8112 9216 8176 9220
rect 8192 9276 8256 9280
rect 8192 9220 8196 9276
rect 8196 9220 8252 9276
rect 8252 9220 8256 9276
rect 8192 9216 8256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 4612 8732 4676 8736
rect 4612 8676 4616 8732
rect 4616 8676 4672 8732
rect 4672 8676 4676 8732
rect 4612 8672 4676 8676
rect 4692 8732 4756 8736
rect 4692 8676 4696 8732
rect 4696 8676 4752 8732
rect 4752 8676 4756 8732
rect 4692 8672 4756 8676
rect 4772 8732 4836 8736
rect 4772 8676 4776 8732
rect 4776 8676 4832 8732
rect 4832 8676 4836 8732
rect 4772 8672 4836 8676
rect 4852 8732 4916 8736
rect 4852 8676 4856 8732
rect 4856 8676 4912 8732
rect 4912 8676 4916 8732
rect 4852 8672 4916 8676
rect 6612 8732 6676 8736
rect 6612 8676 6616 8732
rect 6616 8676 6672 8732
rect 6672 8676 6676 8732
rect 6612 8672 6676 8676
rect 6692 8732 6756 8736
rect 6692 8676 6696 8732
rect 6696 8676 6752 8732
rect 6752 8676 6756 8732
rect 6692 8672 6756 8676
rect 6772 8732 6836 8736
rect 6772 8676 6776 8732
rect 6776 8676 6832 8732
rect 6832 8676 6836 8732
rect 6772 8672 6836 8676
rect 6852 8732 6916 8736
rect 6852 8676 6856 8732
rect 6856 8676 6912 8732
rect 6912 8676 6916 8732
rect 6852 8672 6916 8676
rect 8612 8732 8676 8736
rect 8612 8676 8616 8732
rect 8616 8676 8672 8732
rect 8672 8676 8676 8732
rect 8612 8672 8676 8676
rect 8692 8732 8756 8736
rect 8692 8676 8696 8732
rect 8696 8676 8752 8732
rect 8752 8676 8756 8732
rect 8692 8672 8756 8676
rect 8772 8732 8836 8736
rect 8772 8676 8776 8732
rect 8776 8676 8832 8732
rect 8832 8676 8836 8732
rect 8772 8672 8836 8676
rect 8852 8732 8916 8736
rect 8852 8676 8856 8732
rect 8856 8676 8912 8732
rect 8912 8676 8916 8732
rect 8852 8672 8916 8676
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 3952 8188 4016 8192
rect 3952 8132 3956 8188
rect 3956 8132 4012 8188
rect 4012 8132 4016 8188
rect 3952 8128 4016 8132
rect 4032 8188 4096 8192
rect 4032 8132 4036 8188
rect 4036 8132 4092 8188
rect 4092 8132 4096 8188
rect 4032 8128 4096 8132
rect 4112 8188 4176 8192
rect 4112 8132 4116 8188
rect 4116 8132 4172 8188
rect 4172 8132 4176 8188
rect 4112 8128 4176 8132
rect 4192 8188 4256 8192
rect 4192 8132 4196 8188
rect 4196 8132 4252 8188
rect 4252 8132 4256 8188
rect 4192 8128 4256 8132
rect 5952 8188 6016 8192
rect 5952 8132 5956 8188
rect 5956 8132 6012 8188
rect 6012 8132 6016 8188
rect 5952 8128 6016 8132
rect 6032 8188 6096 8192
rect 6032 8132 6036 8188
rect 6036 8132 6092 8188
rect 6092 8132 6096 8188
rect 6032 8128 6096 8132
rect 6112 8188 6176 8192
rect 6112 8132 6116 8188
rect 6116 8132 6172 8188
rect 6172 8132 6176 8188
rect 6112 8128 6176 8132
rect 6192 8188 6256 8192
rect 6192 8132 6196 8188
rect 6196 8132 6252 8188
rect 6252 8132 6256 8188
rect 6192 8128 6256 8132
rect 7952 8188 8016 8192
rect 7952 8132 7956 8188
rect 7956 8132 8012 8188
rect 8012 8132 8016 8188
rect 7952 8128 8016 8132
rect 8032 8188 8096 8192
rect 8032 8132 8036 8188
rect 8036 8132 8092 8188
rect 8092 8132 8096 8188
rect 8032 8128 8096 8132
rect 8112 8188 8176 8192
rect 8112 8132 8116 8188
rect 8116 8132 8172 8188
rect 8172 8132 8176 8188
rect 8112 8128 8176 8132
rect 8192 8188 8256 8192
rect 8192 8132 8196 8188
rect 8196 8132 8252 8188
rect 8252 8132 8256 8188
rect 8192 8128 8256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 4612 7644 4676 7648
rect 4612 7588 4616 7644
rect 4616 7588 4672 7644
rect 4672 7588 4676 7644
rect 4612 7584 4676 7588
rect 4692 7644 4756 7648
rect 4692 7588 4696 7644
rect 4696 7588 4752 7644
rect 4752 7588 4756 7644
rect 4692 7584 4756 7588
rect 4772 7644 4836 7648
rect 4772 7588 4776 7644
rect 4776 7588 4832 7644
rect 4832 7588 4836 7644
rect 4772 7584 4836 7588
rect 4852 7644 4916 7648
rect 4852 7588 4856 7644
rect 4856 7588 4912 7644
rect 4912 7588 4916 7644
rect 4852 7584 4916 7588
rect 6612 7644 6676 7648
rect 6612 7588 6616 7644
rect 6616 7588 6672 7644
rect 6672 7588 6676 7644
rect 6612 7584 6676 7588
rect 6692 7644 6756 7648
rect 6692 7588 6696 7644
rect 6696 7588 6752 7644
rect 6752 7588 6756 7644
rect 6692 7584 6756 7588
rect 6772 7644 6836 7648
rect 6772 7588 6776 7644
rect 6776 7588 6832 7644
rect 6832 7588 6836 7644
rect 6772 7584 6836 7588
rect 6852 7644 6916 7648
rect 6852 7588 6856 7644
rect 6856 7588 6912 7644
rect 6912 7588 6916 7644
rect 6852 7584 6916 7588
rect 8612 7644 8676 7648
rect 8612 7588 8616 7644
rect 8616 7588 8672 7644
rect 8672 7588 8676 7644
rect 8612 7584 8676 7588
rect 8692 7644 8756 7648
rect 8692 7588 8696 7644
rect 8696 7588 8752 7644
rect 8752 7588 8756 7644
rect 8692 7584 8756 7588
rect 8772 7644 8836 7648
rect 8772 7588 8776 7644
rect 8776 7588 8832 7644
rect 8832 7588 8836 7644
rect 8772 7584 8836 7588
rect 8852 7644 8916 7648
rect 8852 7588 8856 7644
rect 8856 7588 8912 7644
rect 8912 7588 8916 7644
rect 8852 7584 8916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 3952 7100 4016 7104
rect 3952 7044 3956 7100
rect 3956 7044 4012 7100
rect 4012 7044 4016 7100
rect 3952 7040 4016 7044
rect 4032 7100 4096 7104
rect 4032 7044 4036 7100
rect 4036 7044 4092 7100
rect 4092 7044 4096 7100
rect 4032 7040 4096 7044
rect 4112 7100 4176 7104
rect 4112 7044 4116 7100
rect 4116 7044 4172 7100
rect 4172 7044 4176 7100
rect 4112 7040 4176 7044
rect 4192 7100 4256 7104
rect 4192 7044 4196 7100
rect 4196 7044 4252 7100
rect 4252 7044 4256 7100
rect 4192 7040 4256 7044
rect 5952 7100 6016 7104
rect 5952 7044 5956 7100
rect 5956 7044 6012 7100
rect 6012 7044 6016 7100
rect 5952 7040 6016 7044
rect 6032 7100 6096 7104
rect 6032 7044 6036 7100
rect 6036 7044 6092 7100
rect 6092 7044 6096 7100
rect 6032 7040 6096 7044
rect 6112 7100 6176 7104
rect 6112 7044 6116 7100
rect 6116 7044 6172 7100
rect 6172 7044 6176 7100
rect 6112 7040 6176 7044
rect 6192 7100 6256 7104
rect 6192 7044 6196 7100
rect 6196 7044 6252 7100
rect 6252 7044 6256 7100
rect 6192 7040 6256 7044
rect 7952 7100 8016 7104
rect 7952 7044 7956 7100
rect 7956 7044 8012 7100
rect 8012 7044 8016 7100
rect 7952 7040 8016 7044
rect 8032 7100 8096 7104
rect 8032 7044 8036 7100
rect 8036 7044 8092 7100
rect 8092 7044 8096 7100
rect 8032 7040 8096 7044
rect 8112 7100 8176 7104
rect 8112 7044 8116 7100
rect 8116 7044 8172 7100
rect 8172 7044 8176 7100
rect 8112 7040 8176 7044
rect 8192 7100 8256 7104
rect 8192 7044 8196 7100
rect 8196 7044 8252 7100
rect 8252 7044 8256 7100
rect 8192 7040 8256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 4612 6556 4676 6560
rect 4612 6500 4616 6556
rect 4616 6500 4672 6556
rect 4672 6500 4676 6556
rect 4612 6496 4676 6500
rect 4692 6556 4756 6560
rect 4692 6500 4696 6556
rect 4696 6500 4752 6556
rect 4752 6500 4756 6556
rect 4692 6496 4756 6500
rect 4772 6556 4836 6560
rect 4772 6500 4776 6556
rect 4776 6500 4832 6556
rect 4832 6500 4836 6556
rect 4772 6496 4836 6500
rect 4852 6556 4916 6560
rect 4852 6500 4856 6556
rect 4856 6500 4912 6556
rect 4912 6500 4916 6556
rect 4852 6496 4916 6500
rect 6612 6556 6676 6560
rect 6612 6500 6616 6556
rect 6616 6500 6672 6556
rect 6672 6500 6676 6556
rect 6612 6496 6676 6500
rect 6692 6556 6756 6560
rect 6692 6500 6696 6556
rect 6696 6500 6752 6556
rect 6752 6500 6756 6556
rect 6692 6496 6756 6500
rect 6772 6556 6836 6560
rect 6772 6500 6776 6556
rect 6776 6500 6832 6556
rect 6832 6500 6836 6556
rect 6772 6496 6836 6500
rect 6852 6556 6916 6560
rect 6852 6500 6856 6556
rect 6856 6500 6912 6556
rect 6912 6500 6916 6556
rect 6852 6496 6916 6500
rect 8612 6556 8676 6560
rect 8612 6500 8616 6556
rect 8616 6500 8672 6556
rect 8672 6500 8676 6556
rect 8612 6496 8676 6500
rect 8692 6556 8756 6560
rect 8692 6500 8696 6556
rect 8696 6500 8752 6556
rect 8752 6500 8756 6556
rect 8692 6496 8756 6500
rect 8772 6556 8836 6560
rect 8772 6500 8776 6556
rect 8776 6500 8832 6556
rect 8832 6500 8836 6556
rect 8772 6496 8836 6500
rect 8852 6556 8916 6560
rect 8852 6500 8856 6556
rect 8856 6500 8912 6556
rect 8912 6500 8916 6556
rect 8852 6496 8916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 3952 6012 4016 6016
rect 3952 5956 3956 6012
rect 3956 5956 4012 6012
rect 4012 5956 4016 6012
rect 3952 5952 4016 5956
rect 4032 6012 4096 6016
rect 4032 5956 4036 6012
rect 4036 5956 4092 6012
rect 4092 5956 4096 6012
rect 4032 5952 4096 5956
rect 4112 6012 4176 6016
rect 4112 5956 4116 6012
rect 4116 5956 4172 6012
rect 4172 5956 4176 6012
rect 4112 5952 4176 5956
rect 4192 6012 4256 6016
rect 4192 5956 4196 6012
rect 4196 5956 4252 6012
rect 4252 5956 4256 6012
rect 4192 5952 4256 5956
rect 5952 6012 6016 6016
rect 5952 5956 5956 6012
rect 5956 5956 6012 6012
rect 6012 5956 6016 6012
rect 5952 5952 6016 5956
rect 6032 6012 6096 6016
rect 6032 5956 6036 6012
rect 6036 5956 6092 6012
rect 6092 5956 6096 6012
rect 6032 5952 6096 5956
rect 6112 6012 6176 6016
rect 6112 5956 6116 6012
rect 6116 5956 6172 6012
rect 6172 5956 6176 6012
rect 6112 5952 6176 5956
rect 6192 6012 6256 6016
rect 6192 5956 6196 6012
rect 6196 5956 6252 6012
rect 6252 5956 6256 6012
rect 6192 5952 6256 5956
rect 7952 6012 8016 6016
rect 7952 5956 7956 6012
rect 7956 5956 8012 6012
rect 8012 5956 8016 6012
rect 7952 5952 8016 5956
rect 8032 6012 8096 6016
rect 8032 5956 8036 6012
rect 8036 5956 8092 6012
rect 8092 5956 8096 6012
rect 8032 5952 8096 5956
rect 8112 6012 8176 6016
rect 8112 5956 8116 6012
rect 8116 5956 8172 6012
rect 8172 5956 8176 6012
rect 8112 5952 8176 5956
rect 8192 6012 8256 6016
rect 8192 5956 8196 6012
rect 8196 5956 8252 6012
rect 8252 5956 8256 6012
rect 8192 5952 8256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 4612 5468 4676 5472
rect 4612 5412 4616 5468
rect 4616 5412 4672 5468
rect 4672 5412 4676 5468
rect 4612 5408 4676 5412
rect 4692 5468 4756 5472
rect 4692 5412 4696 5468
rect 4696 5412 4752 5468
rect 4752 5412 4756 5468
rect 4692 5408 4756 5412
rect 4772 5468 4836 5472
rect 4772 5412 4776 5468
rect 4776 5412 4832 5468
rect 4832 5412 4836 5468
rect 4772 5408 4836 5412
rect 4852 5468 4916 5472
rect 4852 5412 4856 5468
rect 4856 5412 4912 5468
rect 4912 5412 4916 5468
rect 4852 5408 4916 5412
rect 6612 5468 6676 5472
rect 6612 5412 6616 5468
rect 6616 5412 6672 5468
rect 6672 5412 6676 5468
rect 6612 5408 6676 5412
rect 6692 5468 6756 5472
rect 6692 5412 6696 5468
rect 6696 5412 6752 5468
rect 6752 5412 6756 5468
rect 6692 5408 6756 5412
rect 6772 5468 6836 5472
rect 6772 5412 6776 5468
rect 6776 5412 6832 5468
rect 6832 5412 6836 5468
rect 6772 5408 6836 5412
rect 6852 5468 6916 5472
rect 6852 5412 6856 5468
rect 6856 5412 6912 5468
rect 6912 5412 6916 5468
rect 6852 5408 6916 5412
rect 8612 5468 8676 5472
rect 8612 5412 8616 5468
rect 8616 5412 8672 5468
rect 8672 5412 8676 5468
rect 8612 5408 8676 5412
rect 8692 5468 8756 5472
rect 8692 5412 8696 5468
rect 8696 5412 8752 5468
rect 8752 5412 8756 5468
rect 8692 5408 8756 5412
rect 8772 5468 8836 5472
rect 8772 5412 8776 5468
rect 8776 5412 8832 5468
rect 8832 5412 8836 5468
rect 8772 5408 8836 5412
rect 8852 5468 8916 5472
rect 8852 5412 8856 5468
rect 8856 5412 8912 5468
rect 8912 5412 8916 5468
rect 8852 5408 8916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 3952 4924 4016 4928
rect 3952 4868 3956 4924
rect 3956 4868 4012 4924
rect 4012 4868 4016 4924
rect 3952 4864 4016 4868
rect 4032 4924 4096 4928
rect 4032 4868 4036 4924
rect 4036 4868 4092 4924
rect 4092 4868 4096 4924
rect 4032 4864 4096 4868
rect 4112 4924 4176 4928
rect 4112 4868 4116 4924
rect 4116 4868 4172 4924
rect 4172 4868 4176 4924
rect 4112 4864 4176 4868
rect 4192 4924 4256 4928
rect 4192 4868 4196 4924
rect 4196 4868 4252 4924
rect 4252 4868 4256 4924
rect 4192 4864 4256 4868
rect 5952 4924 6016 4928
rect 5952 4868 5956 4924
rect 5956 4868 6012 4924
rect 6012 4868 6016 4924
rect 5952 4864 6016 4868
rect 6032 4924 6096 4928
rect 6032 4868 6036 4924
rect 6036 4868 6092 4924
rect 6092 4868 6096 4924
rect 6032 4864 6096 4868
rect 6112 4924 6176 4928
rect 6112 4868 6116 4924
rect 6116 4868 6172 4924
rect 6172 4868 6176 4924
rect 6112 4864 6176 4868
rect 6192 4924 6256 4928
rect 6192 4868 6196 4924
rect 6196 4868 6252 4924
rect 6252 4868 6256 4924
rect 6192 4864 6256 4868
rect 7952 4924 8016 4928
rect 7952 4868 7956 4924
rect 7956 4868 8012 4924
rect 8012 4868 8016 4924
rect 7952 4864 8016 4868
rect 8032 4924 8096 4928
rect 8032 4868 8036 4924
rect 8036 4868 8092 4924
rect 8092 4868 8096 4924
rect 8032 4864 8096 4868
rect 8112 4924 8176 4928
rect 8112 4868 8116 4924
rect 8116 4868 8172 4924
rect 8172 4868 8176 4924
rect 8112 4864 8176 4868
rect 8192 4924 8256 4928
rect 8192 4868 8196 4924
rect 8196 4868 8252 4924
rect 8252 4868 8256 4924
rect 8192 4864 8256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 4612 4380 4676 4384
rect 4612 4324 4616 4380
rect 4616 4324 4672 4380
rect 4672 4324 4676 4380
rect 4612 4320 4676 4324
rect 4692 4380 4756 4384
rect 4692 4324 4696 4380
rect 4696 4324 4752 4380
rect 4752 4324 4756 4380
rect 4692 4320 4756 4324
rect 4772 4380 4836 4384
rect 4772 4324 4776 4380
rect 4776 4324 4832 4380
rect 4832 4324 4836 4380
rect 4772 4320 4836 4324
rect 4852 4380 4916 4384
rect 4852 4324 4856 4380
rect 4856 4324 4912 4380
rect 4912 4324 4916 4380
rect 4852 4320 4916 4324
rect 6612 4380 6676 4384
rect 6612 4324 6616 4380
rect 6616 4324 6672 4380
rect 6672 4324 6676 4380
rect 6612 4320 6676 4324
rect 6692 4380 6756 4384
rect 6692 4324 6696 4380
rect 6696 4324 6752 4380
rect 6752 4324 6756 4380
rect 6692 4320 6756 4324
rect 6772 4380 6836 4384
rect 6772 4324 6776 4380
rect 6776 4324 6832 4380
rect 6832 4324 6836 4380
rect 6772 4320 6836 4324
rect 6852 4380 6916 4384
rect 6852 4324 6856 4380
rect 6856 4324 6912 4380
rect 6912 4324 6916 4380
rect 6852 4320 6916 4324
rect 8612 4380 8676 4384
rect 8612 4324 8616 4380
rect 8616 4324 8672 4380
rect 8672 4324 8676 4380
rect 8612 4320 8676 4324
rect 8692 4380 8756 4384
rect 8692 4324 8696 4380
rect 8696 4324 8752 4380
rect 8752 4324 8756 4380
rect 8692 4320 8756 4324
rect 8772 4380 8836 4384
rect 8772 4324 8776 4380
rect 8776 4324 8832 4380
rect 8832 4324 8836 4380
rect 8772 4320 8836 4324
rect 8852 4380 8916 4384
rect 8852 4324 8856 4380
rect 8856 4324 8912 4380
rect 8912 4324 8916 4380
rect 8852 4320 8916 4324
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 3952 3836 4016 3840
rect 3952 3780 3956 3836
rect 3956 3780 4012 3836
rect 4012 3780 4016 3836
rect 3952 3776 4016 3780
rect 4032 3836 4096 3840
rect 4032 3780 4036 3836
rect 4036 3780 4092 3836
rect 4092 3780 4096 3836
rect 4032 3776 4096 3780
rect 4112 3836 4176 3840
rect 4112 3780 4116 3836
rect 4116 3780 4172 3836
rect 4172 3780 4176 3836
rect 4112 3776 4176 3780
rect 4192 3836 4256 3840
rect 4192 3780 4196 3836
rect 4196 3780 4252 3836
rect 4252 3780 4256 3836
rect 4192 3776 4256 3780
rect 5952 3836 6016 3840
rect 5952 3780 5956 3836
rect 5956 3780 6012 3836
rect 6012 3780 6016 3836
rect 5952 3776 6016 3780
rect 6032 3836 6096 3840
rect 6032 3780 6036 3836
rect 6036 3780 6092 3836
rect 6092 3780 6096 3836
rect 6032 3776 6096 3780
rect 6112 3836 6176 3840
rect 6112 3780 6116 3836
rect 6116 3780 6172 3836
rect 6172 3780 6176 3836
rect 6112 3776 6176 3780
rect 6192 3836 6256 3840
rect 6192 3780 6196 3836
rect 6196 3780 6252 3836
rect 6252 3780 6256 3836
rect 6192 3776 6256 3780
rect 7952 3836 8016 3840
rect 7952 3780 7956 3836
rect 7956 3780 8012 3836
rect 8012 3780 8016 3836
rect 7952 3776 8016 3780
rect 8032 3836 8096 3840
rect 8032 3780 8036 3836
rect 8036 3780 8092 3836
rect 8092 3780 8096 3836
rect 8032 3776 8096 3780
rect 8112 3836 8176 3840
rect 8112 3780 8116 3836
rect 8116 3780 8172 3836
rect 8172 3780 8176 3836
rect 8112 3776 8176 3780
rect 8192 3836 8256 3840
rect 8192 3780 8196 3836
rect 8196 3780 8252 3836
rect 8252 3780 8256 3836
rect 8192 3776 8256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 4612 3292 4676 3296
rect 4612 3236 4616 3292
rect 4616 3236 4672 3292
rect 4672 3236 4676 3292
rect 4612 3232 4676 3236
rect 4692 3292 4756 3296
rect 4692 3236 4696 3292
rect 4696 3236 4752 3292
rect 4752 3236 4756 3292
rect 4692 3232 4756 3236
rect 4772 3292 4836 3296
rect 4772 3236 4776 3292
rect 4776 3236 4832 3292
rect 4832 3236 4836 3292
rect 4772 3232 4836 3236
rect 4852 3292 4916 3296
rect 4852 3236 4856 3292
rect 4856 3236 4912 3292
rect 4912 3236 4916 3292
rect 4852 3232 4916 3236
rect 6612 3292 6676 3296
rect 6612 3236 6616 3292
rect 6616 3236 6672 3292
rect 6672 3236 6676 3292
rect 6612 3232 6676 3236
rect 6692 3292 6756 3296
rect 6692 3236 6696 3292
rect 6696 3236 6752 3292
rect 6752 3236 6756 3292
rect 6692 3232 6756 3236
rect 6772 3292 6836 3296
rect 6772 3236 6776 3292
rect 6776 3236 6832 3292
rect 6832 3236 6836 3292
rect 6772 3232 6836 3236
rect 6852 3292 6916 3296
rect 6852 3236 6856 3292
rect 6856 3236 6912 3292
rect 6912 3236 6916 3292
rect 6852 3232 6916 3236
rect 8612 3292 8676 3296
rect 8612 3236 8616 3292
rect 8616 3236 8672 3292
rect 8672 3236 8676 3292
rect 8612 3232 8676 3236
rect 8692 3292 8756 3296
rect 8692 3236 8696 3292
rect 8696 3236 8752 3292
rect 8752 3236 8756 3292
rect 8692 3232 8756 3236
rect 8772 3292 8836 3296
rect 8772 3236 8776 3292
rect 8776 3236 8832 3292
rect 8832 3236 8836 3292
rect 8772 3232 8836 3236
rect 8852 3292 8916 3296
rect 8852 3236 8856 3292
rect 8856 3236 8912 3292
rect 8912 3236 8916 3292
rect 8852 3232 8916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 3952 2748 4016 2752
rect 3952 2692 3956 2748
rect 3956 2692 4012 2748
rect 4012 2692 4016 2748
rect 3952 2688 4016 2692
rect 4032 2748 4096 2752
rect 4032 2692 4036 2748
rect 4036 2692 4092 2748
rect 4092 2692 4096 2748
rect 4032 2688 4096 2692
rect 4112 2748 4176 2752
rect 4112 2692 4116 2748
rect 4116 2692 4172 2748
rect 4172 2692 4176 2748
rect 4112 2688 4176 2692
rect 4192 2748 4256 2752
rect 4192 2692 4196 2748
rect 4196 2692 4252 2748
rect 4252 2692 4256 2748
rect 4192 2688 4256 2692
rect 5952 2748 6016 2752
rect 5952 2692 5956 2748
rect 5956 2692 6012 2748
rect 6012 2692 6016 2748
rect 5952 2688 6016 2692
rect 6032 2748 6096 2752
rect 6032 2692 6036 2748
rect 6036 2692 6092 2748
rect 6092 2692 6096 2748
rect 6032 2688 6096 2692
rect 6112 2748 6176 2752
rect 6112 2692 6116 2748
rect 6116 2692 6172 2748
rect 6172 2692 6176 2748
rect 6112 2688 6176 2692
rect 6192 2748 6256 2752
rect 6192 2692 6196 2748
rect 6196 2692 6252 2748
rect 6252 2692 6256 2748
rect 6192 2688 6256 2692
rect 7952 2748 8016 2752
rect 7952 2692 7956 2748
rect 7956 2692 8012 2748
rect 8012 2692 8016 2748
rect 7952 2688 8016 2692
rect 8032 2748 8096 2752
rect 8032 2692 8036 2748
rect 8036 2692 8092 2748
rect 8092 2692 8096 2748
rect 8032 2688 8096 2692
rect 8112 2748 8176 2752
rect 8112 2692 8116 2748
rect 8116 2692 8172 2748
rect 8172 2692 8176 2748
rect 8112 2688 8176 2692
rect 8192 2748 8256 2752
rect 8192 2692 8196 2748
rect 8196 2692 8252 2748
rect 8252 2692 8256 2748
rect 8192 2688 8256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
rect 4612 2204 4676 2208
rect 4612 2148 4616 2204
rect 4616 2148 4672 2204
rect 4672 2148 4676 2204
rect 4612 2144 4676 2148
rect 4692 2204 4756 2208
rect 4692 2148 4696 2204
rect 4696 2148 4752 2204
rect 4752 2148 4756 2204
rect 4692 2144 4756 2148
rect 4772 2204 4836 2208
rect 4772 2148 4776 2204
rect 4776 2148 4832 2204
rect 4832 2148 4836 2204
rect 4772 2144 4836 2148
rect 4852 2204 4916 2208
rect 4852 2148 4856 2204
rect 4856 2148 4912 2204
rect 4912 2148 4916 2204
rect 4852 2144 4916 2148
rect 6612 2204 6676 2208
rect 6612 2148 6616 2204
rect 6616 2148 6672 2204
rect 6672 2148 6676 2204
rect 6612 2144 6676 2148
rect 6692 2204 6756 2208
rect 6692 2148 6696 2204
rect 6696 2148 6752 2204
rect 6752 2148 6756 2204
rect 6692 2144 6756 2148
rect 6772 2204 6836 2208
rect 6772 2148 6776 2204
rect 6776 2148 6832 2204
rect 6832 2148 6836 2204
rect 6772 2144 6836 2148
rect 6852 2204 6916 2208
rect 6852 2148 6856 2204
rect 6856 2148 6912 2204
rect 6912 2148 6916 2204
rect 6852 2144 6916 2148
rect 8612 2204 8676 2208
rect 8612 2148 8616 2204
rect 8616 2148 8672 2204
rect 8672 2148 8676 2204
rect 8612 2144 8676 2148
rect 8692 2204 8756 2208
rect 8692 2148 8696 2204
rect 8696 2148 8752 2204
rect 8752 2148 8756 2204
rect 8692 2144 8756 2148
rect 8772 2204 8836 2208
rect 8772 2148 8776 2204
rect 8776 2148 8832 2204
rect 8832 2148 8836 2204
rect 8772 2144 8836 2148
rect 8852 2204 8916 2208
rect 8852 2148 8856 2204
rect 8856 2148 8912 2204
rect 8912 2148 8916 2204
rect 8852 2144 8916 2148
<< metal4 >>
rect 1944 9280 2264 9840
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8958 2264 9216
rect 1944 8722 1986 8958
rect 2222 8722 2264 8958
rect 1944 8192 2264 8722
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7054 2032 7104
rect 2096 7054 2112 7104
rect 2176 7054 2192 7104
rect 2256 7040 2264 7104
rect 1944 6818 1986 7040
rect 2222 6818 2264 7040
rect 1944 6016 2264 6818
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 5150 2264 5952
rect 1944 4928 1986 5150
rect 2222 4928 2264 5150
rect 1944 4864 1952 4928
rect 2016 4864 2032 4914
rect 2096 4864 2112 4914
rect 2176 4864 2192 4914
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 3246 2264 3776
rect 1944 3010 1986 3246
rect 2222 3010 2264 3246
rect 1944 2752 2264 3010
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 9824 2924 9840
rect 2604 9760 2612 9824
rect 2676 9760 2692 9824
rect 2756 9760 2772 9824
rect 2836 9760 2852 9824
rect 2916 9760 2924 9824
rect 2604 9618 2924 9760
rect 2604 9382 2646 9618
rect 2882 9382 2924 9618
rect 2604 8736 2924 9382
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7714 2924 8672
rect 2604 7648 2646 7714
rect 2882 7648 2924 7714
rect 2604 7584 2612 7648
rect 2916 7584 2924 7648
rect 2604 7478 2646 7584
rect 2882 7478 2924 7584
rect 2604 6560 2924 7478
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5810 2924 6496
rect 2604 5574 2646 5810
rect 2882 5574 2924 5810
rect 2604 5472 2924 5574
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3906 2924 4320
rect 2604 3670 2646 3906
rect 2882 3670 2924 3906
rect 2604 3296 2924 3670
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
rect 3944 9280 4264 9840
rect 3944 9216 3952 9280
rect 4016 9216 4032 9280
rect 4096 9216 4112 9280
rect 4176 9216 4192 9280
rect 4256 9216 4264 9280
rect 3944 8958 4264 9216
rect 3944 8722 3986 8958
rect 4222 8722 4264 8958
rect 3944 8192 4264 8722
rect 3944 8128 3952 8192
rect 4016 8128 4032 8192
rect 4096 8128 4112 8192
rect 4176 8128 4192 8192
rect 4256 8128 4264 8192
rect 3944 7104 4264 8128
rect 3944 7040 3952 7104
rect 4016 7054 4032 7104
rect 4096 7054 4112 7104
rect 4176 7054 4192 7104
rect 4256 7040 4264 7104
rect 3944 6818 3986 7040
rect 4222 6818 4264 7040
rect 3944 6016 4264 6818
rect 3944 5952 3952 6016
rect 4016 5952 4032 6016
rect 4096 5952 4112 6016
rect 4176 5952 4192 6016
rect 4256 5952 4264 6016
rect 3944 5150 4264 5952
rect 3944 4928 3986 5150
rect 4222 4928 4264 5150
rect 3944 4864 3952 4928
rect 4016 4864 4032 4914
rect 4096 4864 4112 4914
rect 4176 4864 4192 4914
rect 4256 4864 4264 4928
rect 3944 3840 4264 4864
rect 3944 3776 3952 3840
rect 4016 3776 4032 3840
rect 4096 3776 4112 3840
rect 4176 3776 4192 3840
rect 4256 3776 4264 3840
rect 3944 3246 4264 3776
rect 3944 3010 3986 3246
rect 4222 3010 4264 3246
rect 3944 2752 4264 3010
rect 3944 2688 3952 2752
rect 4016 2688 4032 2752
rect 4096 2688 4112 2752
rect 4176 2688 4192 2752
rect 4256 2688 4264 2752
rect 3944 2128 4264 2688
rect 4604 9824 4924 9840
rect 4604 9760 4612 9824
rect 4676 9760 4692 9824
rect 4756 9760 4772 9824
rect 4836 9760 4852 9824
rect 4916 9760 4924 9824
rect 4604 9618 4924 9760
rect 4604 9382 4646 9618
rect 4882 9382 4924 9618
rect 4604 8736 4924 9382
rect 4604 8672 4612 8736
rect 4676 8672 4692 8736
rect 4756 8672 4772 8736
rect 4836 8672 4852 8736
rect 4916 8672 4924 8736
rect 4604 7714 4924 8672
rect 4604 7648 4646 7714
rect 4882 7648 4924 7714
rect 4604 7584 4612 7648
rect 4916 7584 4924 7648
rect 4604 7478 4646 7584
rect 4882 7478 4924 7584
rect 4604 6560 4924 7478
rect 4604 6496 4612 6560
rect 4676 6496 4692 6560
rect 4756 6496 4772 6560
rect 4836 6496 4852 6560
rect 4916 6496 4924 6560
rect 4604 5810 4924 6496
rect 4604 5574 4646 5810
rect 4882 5574 4924 5810
rect 4604 5472 4924 5574
rect 4604 5408 4612 5472
rect 4676 5408 4692 5472
rect 4756 5408 4772 5472
rect 4836 5408 4852 5472
rect 4916 5408 4924 5472
rect 4604 4384 4924 5408
rect 4604 4320 4612 4384
rect 4676 4320 4692 4384
rect 4756 4320 4772 4384
rect 4836 4320 4852 4384
rect 4916 4320 4924 4384
rect 4604 3906 4924 4320
rect 4604 3670 4646 3906
rect 4882 3670 4924 3906
rect 4604 3296 4924 3670
rect 4604 3232 4612 3296
rect 4676 3232 4692 3296
rect 4756 3232 4772 3296
rect 4836 3232 4852 3296
rect 4916 3232 4924 3296
rect 4604 2208 4924 3232
rect 4604 2144 4612 2208
rect 4676 2144 4692 2208
rect 4756 2144 4772 2208
rect 4836 2144 4852 2208
rect 4916 2144 4924 2208
rect 4604 2128 4924 2144
rect 5944 9280 6264 9840
rect 5944 9216 5952 9280
rect 6016 9216 6032 9280
rect 6096 9216 6112 9280
rect 6176 9216 6192 9280
rect 6256 9216 6264 9280
rect 5944 8958 6264 9216
rect 5944 8722 5986 8958
rect 6222 8722 6264 8958
rect 5944 8192 6264 8722
rect 5944 8128 5952 8192
rect 6016 8128 6032 8192
rect 6096 8128 6112 8192
rect 6176 8128 6192 8192
rect 6256 8128 6264 8192
rect 5944 7104 6264 8128
rect 5944 7040 5952 7104
rect 6016 7054 6032 7104
rect 6096 7054 6112 7104
rect 6176 7054 6192 7104
rect 6256 7040 6264 7104
rect 5944 6818 5986 7040
rect 6222 6818 6264 7040
rect 5944 6016 6264 6818
rect 5944 5952 5952 6016
rect 6016 5952 6032 6016
rect 6096 5952 6112 6016
rect 6176 5952 6192 6016
rect 6256 5952 6264 6016
rect 5944 5150 6264 5952
rect 5944 4928 5986 5150
rect 6222 4928 6264 5150
rect 5944 4864 5952 4928
rect 6016 4864 6032 4914
rect 6096 4864 6112 4914
rect 6176 4864 6192 4914
rect 6256 4864 6264 4928
rect 5944 3840 6264 4864
rect 5944 3776 5952 3840
rect 6016 3776 6032 3840
rect 6096 3776 6112 3840
rect 6176 3776 6192 3840
rect 6256 3776 6264 3840
rect 5944 3246 6264 3776
rect 5944 3010 5986 3246
rect 6222 3010 6264 3246
rect 5944 2752 6264 3010
rect 5944 2688 5952 2752
rect 6016 2688 6032 2752
rect 6096 2688 6112 2752
rect 6176 2688 6192 2752
rect 6256 2688 6264 2752
rect 5944 2128 6264 2688
rect 6604 9824 6924 9840
rect 6604 9760 6612 9824
rect 6676 9760 6692 9824
rect 6756 9760 6772 9824
rect 6836 9760 6852 9824
rect 6916 9760 6924 9824
rect 6604 9618 6924 9760
rect 6604 9382 6646 9618
rect 6882 9382 6924 9618
rect 6604 8736 6924 9382
rect 6604 8672 6612 8736
rect 6676 8672 6692 8736
rect 6756 8672 6772 8736
rect 6836 8672 6852 8736
rect 6916 8672 6924 8736
rect 6604 7714 6924 8672
rect 6604 7648 6646 7714
rect 6882 7648 6924 7714
rect 6604 7584 6612 7648
rect 6916 7584 6924 7648
rect 6604 7478 6646 7584
rect 6882 7478 6924 7584
rect 6604 6560 6924 7478
rect 6604 6496 6612 6560
rect 6676 6496 6692 6560
rect 6756 6496 6772 6560
rect 6836 6496 6852 6560
rect 6916 6496 6924 6560
rect 6604 5810 6924 6496
rect 6604 5574 6646 5810
rect 6882 5574 6924 5810
rect 6604 5472 6924 5574
rect 6604 5408 6612 5472
rect 6676 5408 6692 5472
rect 6756 5408 6772 5472
rect 6836 5408 6852 5472
rect 6916 5408 6924 5472
rect 6604 4384 6924 5408
rect 6604 4320 6612 4384
rect 6676 4320 6692 4384
rect 6756 4320 6772 4384
rect 6836 4320 6852 4384
rect 6916 4320 6924 4384
rect 6604 3906 6924 4320
rect 6604 3670 6646 3906
rect 6882 3670 6924 3906
rect 6604 3296 6924 3670
rect 6604 3232 6612 3296
rect 6676 3232 6692 3296
rect 6756 3232 6772 3296
rect 6836 3232 6852 3296
rect 6916 3232 6924 3296
rect 6604 2208 6924 3232
rect 6604 2144 6612 2208
rect 6676 2144 6692 2208
rect 6756 2144 6772 2208
rect 6836 2144 6852 2208
rect 6916 2144 6924 2208
rect 6604 2128 6924 2144
rect 7944 9280 8264 9840
rect 7944 9216 7952 9280
rect 8016 9216 8032 9280
rect 8096 9216 8112 9280
rect 8176 9216 8192 9280
rect 8256 9216 8264 9280
rect 7944 8958 8264 9216
rect 7944 8722 7986 8958
rect 8222 8722 8264 8958
rect 7944 8192 8264 8722
rect 7944 8128 7952 8192
rect 8016 8128 8032 8192
rect 8096 8128 8112 8192
rect 8176 8128 8192 8192
rect 8256 8128 8264 8192
rect 7944 7104 8264 8128
rect 7944 7040 7952 7104
rect 8016 7054 8032 7104
rect 8096 7054 8112 7104
rect 8176 7054 8192 7104
rect 8256 7040 8264 7104
rect 7944 6818 7986 7040
rect 8222 6818 8264 7040
rect 7944 6016 8264 6818
rect 7944 5952 7952 6016
rect 8016 5952 8032 6016
rect 8096 5952 8112 6016
rect 8176 5952 8192 6016
rect 8256 5952 8264 6016
rect 7944 5150 8264 5952
rect 7944 4928 7986 5150
rect 8222 4928 8264 5150
rect 7944 4864 7952 4928
rect 8016 4864 8032 4914
rect 8096 4864 8112 4914
rect 8176 4864 8192 4914
rect 8256 4864 8264 4928
rect 7944 3840 8264 4864
rect 7944 3776 7952 3840
rect 8016 3776 8032 3840
rect 8096 3776 8112 3840
rect 8176 3776 8192 3840
rect 8256 3776 8264 3840
rect 7944 3246 8264 3776
rect 7944 3010 7986 3246
rect 8222 3010 8264 3246
rect 7944 2752 8264 3010
rect 7944 2688 7952 2752
rect 8016 2688 8032 2752
rect 8096 2688 8112 2752
rect 8176 2688 8192 2752
rect 8256 2688 8264 2752
rect 7944 2128 8264 2688
rect 8604 9824 8924 9840
rect 8604 9760 8612 9824
rect 8676 9760 8692 9824
rect 8756 9760 8772 9824
rect 8836 9760 8852 9824
rect 8916 9760 8924 9824
rect 8604 9618 8924 9760
rect 8604 9382 8646 9618
rect 8882 9382 8924 9618
rect 8604 8736 8924 9382
rect 8604 8672 8612 8736
rect 8676 8672 8692 8736
rect 8756 8672 8772 8736
rect 8836 8672 8852 8736
rect 8916 8672 8924 8736
rect 8604 7714 8924 8672
rect 8604 7648 8646 7714
rect 8882 7648 8924 7714
rect 8604 7584 8612 7648
rect 8916 7584 8924 7648
rect 8604 7478 8646 7584
rect 8882 7478 8924 7584
rect 8604 6560 8924 7478
rect 8604 6496 8612 6560
rect 8676 6496 8692 6560
rect 8756 6496 8772 6560
rect 8836 6496 8852 6560
rect 8916 6496 8924 6560
rect 8604 5810 8924 6496
rect 8604 5574 8646 5810
rect 8882 5574 8924 5810
rect 8604 5472 8924 5574
rect 8604 5408 8612 5472
rect 8676 5408 8692 5472
rect 8756 5408 8772 5472
rect 8836 5408 8852 5472
rect 8916 5408 8924 5472
rect 8604 4384 8924 5408
rect 8604 4320 8612 4384
rect 8676 4320 8692 4384
rect 8756 4320 8772 4384
rect 8836 4320 8852 4384
rect 8916 4320 8924 4384
rect 8604 3906 8924 4320
rect 8604 3670 8646 3906
rect 8882 3670 8924 3906
rect 8604 3296 8924 3670
rect 8604 3232 8612 3296
rect 8676 3232 8692 3296
rect 8756 3232 8772 3296
rect 8836 3232 8852 3296
rect 8916 3232 8924 3296
rect 8604 2208 8924 3232
rect 8604 2144 8612 2208
rect 8676 2144 8692 2208
rect 8756 2144 8772 2208
rect 8836 2144 8852 2208
rect 8916 2144 8924 2208
rect 8604 2128 8924 2144
<< via4 >>
rect 1986 8722 2222 8958
rect 1986 7040 2016 7054
rect 2016 7040 2032 7054
rect 2032 7040 2096 7054
rect 2096 7040 2112 7054
rect 2112 7040 2176 7054
rect 2176 7040 2192 7054
rect 2192 7040 2222 7054
rect 1986 6818 2222 7040
rect 1986 4928 2222 5150
rect 1986 4914 2016 4928
rect 2016 4914 2032 4928
rect 2032 4914 2096 4928
rect 2096 4914 2112 4928
rect 2112 4914 2176 4928
rect 2176 4914 2192 4928
rect 2192 4914 2222 4928
rect 1986 3010 2222 3246
rect 2646 9382 2882 9618
rect 2646 7648 2882 7714
rect 2646 7584 2676 7648
rect 2676 7584 2692 7648
rect 2692 7584 2756 7648
rect 2756 7584 2772 7648
rect 2772 7584 2836 7648
rect 2836 7584 2852 7648
rect 2852 7584 2882 7648
rect 2646 7478 2882 7584
rect 2646 5574 2882 5810
rect 2646 3670 2882 3906
rect 3986 8722 4222 8958
rect 3986 7040 4016 7054
rect 4016 7040 4032 7054
rect 4032 7040 4096 7054
rect 4096 7040 4112 7054
rect 4112 7040 4176 7054
rect 4176 7040 4192 7054
rect 4192 7040 4222 7054
rect 3986 6818 4222 7040
rect 3986 4928 4222 5150
rect 3986 4914 4016 4928
rect 4016 4914 4032 4928
rect 4032 4914 4096 4928
rect 4096 4914 4112 4928
rect 4112 4914 4176 4928
rect 4176 4914 4192 4928
rect 4192 4914 4222 4928
rect 3986 3010 4222 3246
rect 4646 9382 4882 9618
rect 4646 7648 4882 7714
rect 4646 7584 4676 7648
rect 4676 7584 4692 7648
rect 4692 7584 4756 7648
rect 4756 7584 4772 7648
rect 4772 7584 4836 7648
rect 4836 7584 4852 7648
rect 4852 7584 4882 7648
rect 4646 7478 4882 7584
rect 4646 5574 4882 5810
rect 4646 3670 4882 3906
rect 5986 8722 6222 8958
rect 5986 7040 6016 7054
rect 6016 7040 6032 7054
rect 6032 7040 6096 7054
rect 6096 7040 6112 7054
rect 6112 7040 6176 7054
rect 6176 7040 6192 7054
rect 6192 7040 6222 7054
rect 5986 6818 6222 7040
rect 5986 4928 6222 5150
rect 5986 4914 6016 4928
rect 6016 4914 6032 4928
rect 6032 4914 6096 4928
rect 6096 4914 6112 4928
rect 6112 4914 6176 4928
rect 6176 4914 6192 4928
rect 6192 4914 6222 4928
rect 5986 3010 6222 3246
rect 6646 9382 6882 9618
rect 6646 7648 6882 7714
rect 6646 7584 6676 7648
rect 6676 7584 6692 7648
rect 6692 7584 6756 7648
rect 6756 7584 6772 7648
rect 6772 7584 6836 7648
rect 6836 7584 6852 7648
rect 6852 7584 6882 7648
rect 6646 7478 6882 7584
rect 6646 5574 6882 5810
rect 6646 3670 6882 3906
rect 7986 8722 8222 8958
rect 7986 7040 8016 7054
rect 8016 7040 8032 7054
rect 8032 7040 8096 7054
rect 8096 7040 8112 7054
rect 8112 7040 8176 7054
rect 8176 7040 8192 7054
rect 8192 7040 8222 7054
rect 7986 6818 8222 7040
rect 7986 4928 8222 5150
rect 7986 4914 8016 4928
rect 8016 4914 8032 4928
rect 8032 4914 8096 4928
rect 8096 4914 8112 4928
rect 8112 4914 8176 4928
rect 8176 4914 8192 4928
rect 8192 4914 8222 4928
rect 7986 3010 8222 3246
rect 8646 9382 8882 9618
rect 8646 7648 8882 7714
rect 8646 7584 8676 7648
rect 8676 7584 8692 7648
rect 8692 7584 8756 7648
rect 8756 7584 8772 7648
rect 8772 7584 8836 7648
rect 8836 7584 8852 7648
rect 8852 7584 8882 7648
rect 8646 7478 8882 7584
rect 8646 5574 8882 5810
rect 8646 3670 8882 3906
<< metal5 >>
rect 1056 9618 9156 9660
rect 1056 9382 2646 9618
rect 2882 9382 4646 9618
rect 4882 9382 6646 9618
rect 6882 9382 8646 9618
rect 8882 9382 9156 9618
rect 1056 9340 9156 9382
rect 1056 8958 9156 9000
rect 1056 8722 1986 8958
rect 2222 8722 3986 8958
rect 4222 8722 5986 8958
rect 6222 8722 7986 8958
rect 8222 8722 9156 8958
rect 1056 8680 9156 8722
rect 1056 7714 9156 7756
rect 1056 7478 2646 7714
rect 2882 7478 4646 7714
rect 4882 7478 6646 7714
rect 6882 7478 8646 7714
rect 8882 7478 9156 7714
rect 1056 7436 9156 7478
rect 1056 7054 9156 7096
rect 1056 6818 1986 7054
rect 2222 6818 3986 7054
rect 4222 6818 5986 7054
rect 6222 6818 7986 7054
rect 8222 6818 9156 7054
rect 1056 6776 9156 6818
rect 1056 5810 9156 5852
rect 1056 5574 2646 5810
rect 2882 5574 4646 5810
rect 4882 5574 6646 5810
rect 6882 5574 8646 5810
rect 8882 5574 9156 5810
rect 1056 5532 9156 5574
rect 1056 5150 9156 5192
rect 1056 4914 1986 5150
rect 2222 4914 3986 5150
rect 4222 4914 5986 5150
rect 6222 4914 7986 5150
rect 8222 4914 9156 5150
rect 1056 4872 9156 4914
rect 1056 3906 9156 3948
rect 1056 3670 2646 3906
rect 2882 3670 4646 3906
rect 4882 3670 6646 3906
rect 6882 3670 8646 3906
rect 8882 3670 9156 3906
rect 1056 3628 9156 3670
rect 1056 3246 9156 3288
rect 1056 3010 1986 3246
rect 2222 3010 3986 3246
rect 4222 3010 5986 3246
rect 6222 3010 7986 3246
rect 8222 3010 9156 3246
rect 1056 2968 9156 3010
use sky130_fd_sc_hd__or3b_2  _053_
timestamp 0
transform 1 0 3036 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _054_
timestamp 0
transform 1 0 5428 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _055_
timestamp 0
transform -1 0 4416 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _056_
timestamp 0
transform 1 0 8372 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _057_
timestamp 0
transform -1 0 8372 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _058_
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _059_
timestamp 0
transform -1 0 4232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _060_
timestamp 0
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _061_
timestamp 0
transform -1 0 5060 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _062_
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _063_
timestamp 0
transform -1 0 7820 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _064_
timestamp 0
transform -1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _065_
timestamp 0
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _066_
timestamp 0
transform -1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _067_
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _068_
timestamp 0
transform 1 0 2576 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _069_
timestamp 0
transform -1 0 5336 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _070_
timestamp 0
transform -1 0 8464 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _071_
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _072_
timestamp 0
transform 1 0 5888 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _073_
timestamp 0
transform 1 0 4416 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _074_
timestamp 0
transform -1 0 5888 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _075_
timestamp 0
transform -1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _076_
timestamp 0
transform 1 0 3036 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _077_
timestamp 0
transform -1 0 3864 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _078_
timestamp 0
transform 1 0 1748 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _079_
timestamp 0
transform -1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _080_
timestamp 0
transform 1 0 2760 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _081_
timestamp 0
transform 1 0 3220 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _082_
timestamp 0
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _083_
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _084_
timestamp 0
transform 1 0 3404 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _085_
timestamp 0
transform -1 0 5888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _086_
timestamp 0
transform 1 0 4600 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _087_
timestamp 0
transform -1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _088_
timestamp 0
transform 1 0 1656 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _089_
timestamp 0
transform 1 0 2024 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _090_
timestamp 0
transform 1 0 4048 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _091_
timestamp 0
transform 1 0 7268 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _092_
timestamp 0
transform 1 0 6348 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _093_
timestamp 0
transform -1 0 8372 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _094_
timestamp 0
transform 1 0 2760 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_1  _095_
timestamp 0
transform 1 0 4784 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _096_
timestamp 0
transform -1 0 6164 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _097_
timestamp 0
transform -1 0 6072 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _098_
timestamp 0
transform 1 0 6072 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _099_
timestamp 0
transform -1 0 7268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _100_
timestamp 0
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _101_
timestamp 0
transform 1 0 6992 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _102_
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _103_
timestamp 0
transform 1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _104_
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _105_
timestamp 0
transform 1 0 4968 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _106_
timestamp 0
transform 1 0 5612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _107_
timestamp 0
transform 1 0 6440 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _108_
timestamp 0
transform 1 0 4048 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 0
transform -1 0 5060 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlxtn_1  _110_
timestamp 0
transform 1 0 5244 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_7
timestamp 0
transform 1 0 1748 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_20
timestamp 0
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49
timestamp 0
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 0
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 0
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_9
timestamp 0
transform 1 0 1932 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_21
timestamp 0
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_52
timestamp 0
transform 1 0 5888 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_64
timestamp 0
transform 1 0 6992 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_57
timestamp 0
transform 1 0 6348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_69
timestamp 0
transform 1 0 7452 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_28
timestamp 0
transform 1 0 3680 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_40
timestamp 0
transform 1 0 4784 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_62
timestamp 0
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_73
timestamp 0
transform 1 0 7820 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_16
timestamp 0
transform 1 0 2576 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_34
timestamp 0
transform 1 0 4232 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_46
timestamp 0
transform 1 0 5336 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_58
timestamp 0
transform 1 0 6440 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_70
timestamp 0
transform 1 0 7544 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_82
timestamp 0
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_9
timestamp 0
transform 1 0 1932 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_24
timestamp 0
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_36
timestamp 0
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_46
timestamp 0
transform 1 0 5336 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 0
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_10
timestamp 0
transform 1 0 2024 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_22
timestamp 0
transform 1 0 3128 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_45
timestamp 0
transform 1 0 5244 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_62
timestamp 0
transform 1 0 6808 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_73
timestamp 0
transform 1 0 7820 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 0
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_22
timestamp 0
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_43
timestamp 0
transform 1 0 5060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_60
timestamp 0
transform 1 0 6624 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_71
timestamp 0
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_79
timestamp 0
transform 1 0 8372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_83
timestamp 0
transform 1 0 8740 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_73
timestamp 0
transform 1 0 7820 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 0
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_22
timestamp 0
transform 1 0 3128 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_34
timestamp 0
transform 1 0 4232 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_46
timestamp 0
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 0
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_63
timestamp 0
transform 1 0 6900 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_75
timestamp 0
transform 1 0 8004 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_16
timestamp 0
transform 1 0 2576 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_37
timestamp 0
transform 1 0 4508 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_52
timestamp 0
transform 1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_56
timestamp 0
transform 1 0 6256 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_72
timestamp 0
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_30
timestamp 0
transform 1 0 3864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_34
timestamp 0
transform 1 0 4232 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_38
timestamp 0
transform 1 0 4600 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_45
timestamp 0
transform 1 0 5244 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 0
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_13
timestamp 0
transform 1 0 2300 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 0
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_43
timestamp 0
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_57
timestamp 0
transform 1 0 6348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_69
timestamp 0
transform 1 0 7452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_81
timestamp 0
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_11
timestamp 0
transform 1 0 2116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_23
timestamp 0
transform 1 0 3220 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_29
timestamp 0
transform 1 0 3772 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_37
timestamp 0
transform 1 0 4508 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 0
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 0
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_65
timestamp 0
transform 1 0 7084 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_72
timestamp 0
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform -1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 0
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 0
transform -1 0 8280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 0
transform -1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform 1 0 4600 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 0
transform 1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 0
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 0
transform 1 0 7176 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 0
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 0
transform -1 0 1932 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 0
transform 1 0 8280 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output16
timestamp 0
transform -1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 9108 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 9108 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 9108 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 9108 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 9108 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 9108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 9108 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 9108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 9108 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 9108 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 9108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 9108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 9108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 0
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
<< labels >>
rlabel metal1 s 5106 9792 5106 9792 4 VGND
rlabel metal1 s 5106 9248 5106 9248 4 VPWR
rlabel metal1 s 5934 3910 5934 3910 4 _000_
rlabel metal1 s 5152 9010 5152 9010 4 _001_
rlabel metal1 s 5796 7854 5796 7854 4 _002_
rlabel metal1 s 5750 3502 5750 3502 4 _003_
rlabel metal1 s 6164 3026 6164 3026 4 _004_
rlabel metal1 s 7774 5780 7774 5780 4 _005_
rlabel metal1 s 6578 6222 6578 6222 4 _006_
rlabel metal1 s 5198 7718 5198 7718 4 _007_
rlabel metal2 s 3726 7276 3726 7276 4 _008_
rlabel metal1 s 4738 6188 4738 6188 4 _009_
rlabel metal1 s 5842 6120 5842 6120 4 _010_
rlabel metal1 s 6624 6086 6624 6086 4 _011_
rlabel metal2 s 7406 4828 7406 4828 4 _012_
rlabel metal1 s 5658 4080 5658 4080 4 _013_
rlabel metal1 s 6118 4080 6118 4080 4 _014_
rlabel metal1 s 6118 6324 6118 6324 4 _015_
rlabel metal1 s 5290 7854 5290 7854 4 _016_
rlabel metal1 s 4094 7514 4094 7514 4 _017_
rlabel metal2 s 6486 7854 6486 7854 4 _018_
rlabel metal1 s 7636 6970 7636 6970 4 _019_
rlabel metal1 s 6440 4182 6440 4182 4 _020_
rlabel metal1 s 5842 3978 5842 3978 4 _021_
rlabel metal1 s 5014 3162 5014 3162 4 _022_
rlabel metal1 s 2254 4556 2254 4556 4 _023_
rlabel metal2 s 3626 8602 3626 8602 4 _024_
rlabel metal2 s 2990 8364 2990 8364 4 _025_
rlabel metal2 s 2162 4318 2162 4318 4 _026_
rlabel metal1 s 3082 8432 3082 8432 4 _027_
rlabel metal1 s 4738 4658 4738 4658 4 _028_
rlabel metal1 s 3274 4454 3274 4454 4 _029_
rlabel metal1 s 5520 5678 5520 5678 4 _030_
rlabel metal1 s 4140 6222 4140 6222 4 _031_
rlabel metal1 s 4830 7412 4830 7412 4 _032_
rlabel metal2 s 4554 6732 4554 6732 4 _033_
rlabel metal1 s 2346 6188 2346 6188 4 _034_
rlabel metal1 s 1886 5542 1886 5542 4 _035_
rlabel metal1 s 4692 6290 4692 6290 4 _036_
rlabel metal1 s 6854 7888 6854 7888 4 _037_
rlabel metal1 s 6762 7888 6762 7888 4 _038_
rlabel metal1 s 6486 5644 6486 5644 4 _039_
rlabel metal1 s 4692 4590 4692 4590 4 _040_
rlabel metal1 s 5704 5338 5704 5338 4 _041_
rlabel metal1 s 5382 5712 5382 5712 4 _042_
rlabel metal1 s 6118 5644 6118 5644 4 _043_
rlabel metal1 s 6900 5882 6900 5882 4 _044_
rlabel metal1 s 7084 2958 7084 2958 4 _045_
rlabel metal1 s 6992 3026 6992 3026 4 _046_
rlabel metal1 s 6463 3502 6463 3502 4 _047_
rlabel metal2 s 4922 4624 4922 4624 4 _048_
rlabel metal1 s 5934 3502 5934 3502 4 _049_
rlabel metal1 s 5520 3162 5520 3162 4 _050_
rlabel metal1 s 6486 3026 6486 3026 4 _051_
rlabel metal1 s 4646 8942 4646 8942 4 _052_
rlabel metal1 s 9016 7378 9016 7378 4 a[0]
rlabel metal3 s 843 11628 843 11628 4 a[1]
rlabel metal1 s 8234 9520 8234 9520 4 a[2]
rlabel metal1 s 8418 2380 8418 2380 4 a[3]
rlabel metal1 s 4600 9554 4600 9554 4 b[0]
rlabel metal2 s 46 1554 46 1554 4 b[1]
rlabel metal2 s 8418 1588 8418 1588 4 b[2]
rlabel metal2 s 2622 1027 2622 1027 4 b[3]
rlabel metal1 s 7544 9622 7544 9622 4 carry
rlabel metal2 s 5014 7752 5014 7752 4 net1
rlabel metal1 s 1656 5882 1656 5882 4 net10
rlabel metal1 s 4186 4046 4186 4046 4 net11
rlabel metal1 s 6808 9146 6808 9146 4 net12
rlabel metal2 s 3174 5712 3174 5712 4 net13
rlabel metal2 s 3450 5678 3450 5678 4 net14
rlabel metal1 s 7498 8058 7498 8058 4 net15
rlabel metal1 s 5980 2414 5980 2414 4 net16
rlabel metal1 s 1702 6324 1702 6324 4 net2
rlabel metal1 s 8050 6868 8050 6868 4 net3
rlabel metal1 s 7728 2618 7728 2618 4 net4
rlabel metal1 s 4876 8466 4876 8466 4 net5
rlabel metal1 s 1702 6426 1702 6426 4 net6
rlabel metal1 s 8602 2618 8602 2618 4 net7
rlabel metal1 s 3542 3026 3542 3026 4 net8
rlabel metal1 s 2392 8942 2392 8942 4 net9
rlabel metal3 s 820 2788 820 2788 4 out[0]
rlabel metal3 s 820 5508 820 5508 4 out[1]
rlabel metal1 s 9246 9622 9246 9622 4 out[2]
rlabel metal2 s 5198 1520 5198 1520 4 out[3]
rlabel metal3 s 820 8908 820 8908 4 sel[0]
rlabel metal1 s 1426 9622 1426 9622 4 sel[1]
rlabel metal1 s 9016 3502 9016 3502 4 sel[2]
flabel metal5 s 1056 9340 9156 9660 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 7436 9156 7756 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 5532 9156 5852 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3628 9156 3948 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 8604 2128 8924 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 6604 2128 6924 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4604 2128 4924 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2604 2128 2924 9840 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 8680 9156 9000 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 6776 9156 7096 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 4872 9156 5192 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 2968 9156 3288 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 7944 2128 8264 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 5944 2128 6264 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 3944 2128 4264 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 1944 2128 2264 9840 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 9474 6808 10274 6928 0 FreeSans 600 0 0 0 a[0]
port 3 nsew
flabel metal3 s 0 11568 800 11688 0 FreeSans 600 0 0 0 a[1]
port 4 nsew
flabel metal3 s 9474 9528 10274 9648 0 FreeSans 600 0 0 0 a[2]
port 5 nsew
flabel metal3 s 9474 688 10274 808 0 FreeSans 600 0 0 0 a[3]
port 6 nsew
flabel metal2 s 4526 11618 4582 12418 0 FreeSans 280 90 0 0 b[0]
port 7 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 b[1]
port 8 nsew
flabel metal2 s 8390 0 8446 800 0 FreeSans 280 90 0 0 b[2]
port 9 nsew
flabel metal2 s 2594 0 2650 800 0 FreeSans 280 90 0 0 b[3]
port 10 nsew
flabel metal2 s 7102 11618 7158 12418 0 FreeSans 280 90 0 0 carry
port 11 nsew
flabel metal3 s 0 2728 800 2848 0 FreeSans 600 0 0 0 out[0]
port 12 nsew
flabel metal3 s 0 5448 800 5568 0 FreeSans 600 0 0 0 out[1]
port 13 nsew
flabel metal2 s 9678 11618 9734 12418 0 FreeSans 280 90 0 0 out[2]
port 14 nsew
flabel metal2 s 5170 0 5226 800 0 FreeSans 280 90 0 0 out[3]
port 15 nsew
flabel metal3 s 0 8848 800 8968 0 FreeSans 600 0 0 0 sel[0]
port 16 nsew
flabel metal2 s 1306 11618 1362 12418 0 FreeSans 280 90 0 0 sel[1]
port 17 nsew
flabel metal3 s 9474 3408 10274 3528 0 FreeSans 600 0 0 0 sel[2]
port 18 nsew
<< properties >>
string FIXED_BBOX 0 0 10274 12418
<< end >>
